------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 3.4
--  \   \         Application : 7 Series FPGAs Transceivers Wizard 
--  /   /         Filename : xlaui_support.vhd
-- /___/   /\      
-- \   \  /  \ 
--  \___\/\___\
--
--  Description : This module instantiates the modules required for
--                reset and initialisation of the Transceiver
--
-- Module XLAUI_support
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;
--***********************************Entity Declaration************************

entity XLAUI_support is
	generic(
		EXAMPLE_SIM_GTRESET_SPEEDUP : string  := "TRUE"; -- simulation setting for GT SecureIP model
		STABLE_CLOCK_PERIOD         : integer := 6
	);
	port(
		--____________________________COMMON PORTS________________________________
		SYS_CLK_I                   : in  std_logic;

		SOFT_RESET_IN               : in  std_logic;
		DONT_RESET_ON_DATA_ERROR_IN : in  std_logic;

		GTREFCLK_PAD_N_IN           : in  std_logic;
		GTREFCLK_PAD_P_IN           : in  std_logic;

		GTREFCLK_O                  : out std_logic;

		GT0_TXOUTCLK_OUT            : out std_logic;
		GT_TXUSRCLK2_IN             : in  std_logic;
		GT_TXUSRCLK_IN              : in  std_logic;
		GT_TXUSRCLK_LOCKED_IN       : in  std_logic;
		GT_TXUSRCLK_RESET_OUT       : out std_logic;

		GT0_RXOUTCLK_OUT            : out std_logic;
		GT_RXUSRCLK2_IN             : in  std_logic;
		GT_RXUSRCLK_IN              : in  std_logic;
		GT_RXUSRCLK_LOCKED_IN       : in  std_logic;
		GT_RXUSRCLK_RESET_OUT       : out std_logic;

		GT0_TX_FSM_RESET_DONE_OUT   : out std_logic;
		GT0_RX_FSM_RESET_DONE_OUT   : out std_logic;
		GT0_DATA_VALID_IN           : in  std_logic;
		GT1_TX_FSM_RESET_DONE_OUT   : out std_logic;
		GT1_RX_FSM_RESET_DONE_OUT   : out std_logic;
		GT1_DATA_VALID_IN           : in  std_logic;
		GT2_TX_FSM_RESET_DONE_OUT   : out std_logic;
		GT2_RX_FSM_RESET_DONE_OUT   : out std_logic;
		GT2_DATA_VALID_IN           : in  std_logic;
		GT3_TX_FSM_RESET_DONE_OUT   : out std_logic;
		GT3_RX_FSM_RESET_DONE_OUT   : out std_logic;
		GT3_DATA_VALID_IN           : in  std_logic;

		--_________________________________________________________________________
		--GT0  (X0Y36)
		--____________________________CHANNEL PORTS________________________________
		---------------------------- Channel - DRP Ports  --------------------------
		gt0_drpaddr_in              : in  std_logic_vector(8 downto 0);
		gt0_drpdi_in                : in  std_logic_vector(15 downto 0);
		gt0_drpdo_out               : out std_logic_vector(15 downto 0);
		gt0_drpen_in                : in  std_logic;
		gt0_drprdy_out              : out std_logic;
		gt0_drpwe_in                : in  std_logic;
		------------------------------- Loopback Ports -----------------------------
		gt0_loopback_in             : in  std_logic_vector(2 downto 0);
		--------------------- RX Initialization and Reset Ports --------------------
		gt0_eyescanreset_in         : in  std_logic;
		gt0_rxuserrdy_in            : in  std_logic;
		-------------------------- RX Margin Analysis Ports ------------------------
		gt0_eyescandataerror_out    : out std_logic;
		gt0_eyescantrigger_in       : in  std_logic;
		------------------- Receive Ports - Digital Monitor Ports ------------------
		gt0_dmonitorout_out         : out std_logic_vector(14 downto 0);
		------------------ Receive Ports - FPGA RX interface Ports -----------------
		gt0_rxdata_out              : out std_logic_vector(63 downto 0);
		------------------- Receive Ports - Pattern Checker Ports ------------------
		gt0_rxprbserr_out           : out std_logic;
		gt0_rxprbssel_in            : in  std_logic_vector(2 downto 0);
		------------------- Receive Ports - Pattern Checker ports ------------------
		gt0_rxprbscntreset_in       : in  std_logic;
		------------------------ Receive Ports - RX AFE Ports ----------------------
		gt0_gthrxn_in               : in  std_logic;
		------------------- Receive Ports - RX Buffer Bypass Ports -----------------
		gt0_rxbufreset_in           : in  std_logic;
		gt0_rxbufstatus_out         : out std_logic_vector(2 downto 0);
		--------------------- Receive Ports - RX Equalizer Ports -------------------
		gt0_rxmonitorout_out        : out std_logic_vector(6 downto 0);
		gt0_rxmonitorsel_in         : in  std_logic_vector(1 downto 0);
		---------------------- Receive Ports - RX Gearbox Ports --------------------
		gt0_rxdatavalid_out         : out std_logic;
		gt0_rxheader_out            : out std_logic_vector(1 downto 0);
		gt0_rxheadervalid_out       : out std_logic;
		--------------------- Receive Ports - RX Gearbox Ports  --------------------
		gt0_rxgearboxslip_in        : in  std_logic;
		------------- Receive Ports - RX Initialization and Reset Ports ------------
		gt0_gtrxreset_in            : in  std_logic;
		gt0_rxpcsreset_in           : in  std_logic;
		------------------------ Receive Ports -RX AFE Ports -----------------------
		gt0_gthrxp_in               : in  std_logic;
		-------------- Receive Ports -RX Initialization and Reset Ports ------------
		gt0_rxresetdone_out         : out std_logic;
		--------------------- TX Initialization and Reset Ports --------------------
		gt0_gttxreset_in            : in  std_logic;
		gt0_txuserrdy_in            : in  std_logic;
		-------------- Transmit Ports - 64b66b and 64b67b Gearbox Ports ------------
		gt0_txheader_in             : in  std_logic_vector(1 downto 0);
		--------------------- Transmit Ports - PCI Express Ports -------------------
		gt0_txelecidle_in           : in  std_logic;
		------------------ Transmit Ports - Pattern Generator Ports ----------------
		gt0_txprbsforceerr_in       : in  std_logic;
		---------------------- Transmit Ports - TX Buffer Ports --------------------
		gt0_txbufstatus_out         : out std_logic_vector(1 downto 0);
		------------------ Transmit Ports - TX Data Path interface -----------------
		gt0_txdata_in               : in  std_logic_vector(63 downto 0);
		---------------- Transmit Ports - TX Driver and OOB signaling --------------
		gt0_gthtxn_out              : out std_logic;
		gt0_gthtxp_out              : out std_logic;
		--------------------- Transmit Ports - TX Gearbox Ports --------------------
		gt0_txsequence_in           : in  std_logic_vector(6 downto 0);
		------------- Transmit Ports - TX Initialization and Reset Ports -----------
		gt0_txpcsreset_in           : in  std_logic;
		gt0_txresetdone_out         : out std_logic;
		----------------- Transmit Ports - TX Polarity Control Ports ---------------
		gt0_txpolarity_in           : in  std_logic;
		------------------ Transmit Ports - pattern Generator Ports ----------------
		gt0_txprbssel_in            : in  std_logic_vector(2 downto 0);

		--GT1  (X0Y37)
		--____________________________CHANNEL PORTS________________________________
		---------------------------- Channel - DRP Ports  --------------------------
		gt1_drpaddr_in              : in  std_logic_vector(8 downto 0);
		gt1_drpdi_in                : in  std_logic_vector(15 downto 0);
		gt1_drpdo_out               : out std_logic_vector(15 downto 0);
		gt1_drpen_in                : in  std_logic;
		gt1_drprdy_out              : out std_logic;
		gt1_drpwe_in                : in  std_logic;
		------------------------------- Loopback Ports -----------------------------
		gt1_loopback_in             : in  std_logic_vector(2 downto 0);
		--------------------- RX Initialization and Reset Ports --------------------
		gt1_eyescanreset_in         : in  std_logic;
		gt1_rxuserrdy_in            : in  std_logic;
		-------------------------- RX Margin Analysis Ports ------------------------
		gt1_eyescandataerror_out    : out std_logic;
		gt1_eyescantrigger_in       : in  std_logic;
		------------------- Receive Ports - Digital Monitor Ports ------------------
		gt1_dmonitorout_out         : out std_logic_vector(14 downto 0);
		------------------ Receive Ports - FPGA RX interface Ports -----------------
		gt1_rxdata_out              : out std_logic_vector(63 downto 0);
		------------------- Receive Ports - Pattern Checker Ports ------------------
		gt1_rxprbserr_out           : out std_logic;
		gt1_rxprbssel_in            : in  std_logic_vector(2 downto 0);
		------------------- Receive Ports - Pattern Checker ports ------------------
		gt1_rxprbscntreset_in       : in  std_logic;
		------------------------ Receive Ports - RX AFE Ports ----------------------
		gt1_gthrxn_in               : in  std_logic;
		------------------- Receive Ports - RX Buffer Bypass Ports -----------------
		gt1_rxbufreset_in           : in  std_logic;
		gt1_rxbufstatus_out         : out std_logic_vector(2 downto 0);
		--------------------- Receive Ports - RX Equalizer Ports -------------------
		gt1_rxmonitorout_out        : out std_logic_vector(6 downto 0);
		gt1_rxmonitorsel_in         : in  std_logic_vector(1 downto 0);
		---------------------- Receive Ports - RX Gearbox Ports --------------------
		gt1_rxdatavalid_out         : out std_logic;
		gt1_rxheader_out            : out std_logic_vector(1 downto 0);
		gt1_rxheadervalid_out       : out std_logic;
		--------------------- Receive Ports - RX Gearbox Ports  --------------------
		gt1_rxgearboxslip_in        : in  std_logic;
		------------- Receive Ports - RX Initialization and Reset Ports ------------
		gt1_gtrxreset_in            : in  std_logic;
		gt1_rxpcsreset_in           : in  std_logic;
		------------------------ Receive Ports -RX AFE Ports -----------------------
		gt1_gthrxp_in               : in  std_logic;
		-------------- Receive Ports -RX Initialization and Reset Ports ------------
		gt1_rxresetdone_out         : out std_logic;
		--------------------- TX Initialization and Reset Ports --------------------
		gt1_gttxreset_in            : in  std_logic;
		gt1_txuserrdy_in            : in  std_logic;
		-------------- Transmit Ports - 64b66b and 64b67b Gearbox Ports ------------
		gt1_txheader_in             : in  std_logic_vector(1 downto 0);
		--------------------- Transmit Ports - PCI Express Ports -------------------
		gt1_txelecidle_in           : in  std_logic;
		------------------ Transmit Ports - Pattern Generator Ports ----------------
		gt1_txprbsforceerr_in       : in  std_logic;
		---------------------- Transmit Ports - TX Buffer Ports --------------------
		gt1_txbufstatus_out         : out std_logic_vector(1 downto 0);
		------------------ Transmit Ports - TX Data Path interface -----------------
		gt1_txdata_in               : in  std_logic_vector(63 downto 0);
		---------------- Transmit Ports - TX Driver and OOB signaling --------------
		gt1_gthtxn_out              : out std_logic;
		gt1_gthtxp_out              : out std_logic;
		--------------------- Transmit Ports - TX Gearbox Ports --------------------
		gt1_txsequence_in           : in  std_logic_vector(6 downto 0);
		------------- Transmit Ports - TX Initialization and Reset Ports -----------
		gt1_txpcsreset_in           : in  std_logic;
		gt1_txresetdone_out         : out std_logic;
		----------------- Transmit Ports - TX Polarity Control Ports ---------------
		gt1_txpolarity_in           : in  std_logic;
		------------------ Transmit Ports - pattern Generator Ports ----------------
		gt1_txprbssel_in            : in  std_logic_vector(2 downto 0);

		--GT2  (X0Y38)
		--____________________________CHANNEL PORTS________________________________
		---------------------------- Channel - DRP Ports  --------------------------
		gt2_drpaddr_in              : in  std_logic_vector(8 downto 0);
		gt2_drpdi_in                : in  std_logic_vector(15 downto 0);
		gt2_drpdo_out               : out std_logic_vector(15 downto 0);
		gt2_drpen_in                : in  std_logic;
		gt2_drprdy_out              : out std_logic;
		gt2_drpwe_in                : in  std_logic;
		------------------------------- Loopback Ports -----------------------------
		gt2_loopback_in             : in  std_logic_vector(2 downto 0);
		--------------------- RX Initialization and Reset Ports --------------------
		gt2_eyescanreset_in         : in  std_logic;
		gt2_rxuserrdy_in            : in  std_logic;
		-------------------------- RX Margin Analysis Ports ------------------------
		gt2_eyescandataerror_out    : out std_logic;
		gt2_eyescantrigger_in       : in  std_logic;
		------------------- Receive Ports - Digital Monitor Ports ------------------
		gt2_dmonitorout_out         : out std_logic_vector(14 downto 0);
		------------------ Receive Ports - FPGA RX interface Ports -----------------
		gt2_rxdata_out              : out std_logic_vector(63 downto 0);
		------------------- Receive Ports - Pattern Checker Ports ------------------
		gt2_rxprbserr_out           : out std_logic;
		gt2_rxprbssel_in            : in  std_logic_vector(2 downto 0);
		------------------- Receive Ports - Pattern Checker ports ------------------
		gt2_rxprbscntreset_in       : in  std_logic;
		------------------------ Receive Ports - RX AFE Ports ----------------------
		gt2_gthrxn_in               : in  std_logic;
		------------------- Receive Ports - RX Buffer Bypass Ports -----------------
		gt2_rxbufreset_in           : in  std_logic;
		gt2_rxbufstatus_out         : out std_logic_vector(2 downto 0);
		--------------------- Receive Ports - RX Equalizer Ports -------------------
		gt2_rxmonitorout_out        : out std_logic_vector(6 downto 0);
		gt2_rxmonitorsel_in         : in  std_logic_vector(1 downto 0);
		---------------------- Receive Ports - RX Gearbox Ports --------------------
		gt2_rxdatavalid_out         : out std_logic;
		gt2_rxheader_out            : out std_logic_vector(1 downto 0);
		gt2_rxheadervalid_out       : out std_logic;
		--------------------- Receive Ports - RX Gearbox Ports  --------------------
		gt2_rxgearboxslip_in        : in  std_logic;
		------------- Receive Ports - RX Initialization and Reset Ports ------------
		gt2_gtrxreset_in            : in  std_logic;
		gt2_rxpcsreset_in           : in  std_logic;
		------------------------ Receive Ports -RX AFE Ports -----------------------
		gt2_gthrxp_in               : in  std_logic;
		-------------- Receive Ports -RX Initialization and Reset Ports ------------
		gt2_rxresetdone_out         : out std_logic;
		--------------------- TX Initialization and Reset Ports --------------------
		gt2_gttxreset_in            : in  std_logic;
		gt2_txuserrdy_in            : in  std_logic;
		-------------- Transmit Ports - 64b66b and 64b67b Gearbox Ports ------------
		gt2_txheader_in             : in  std_logic_vector(1 downto 0);
		--------------------- Transmit Ports - PCI Express Ports -------------------
		gt2_txelecidle_in           : in  std_logic;
		------------------ Transmit Ports - Pattern Generator Ports ----------------
		gt2_txprbsforceerr_in       : in  std_logic;
		---------------------- Transmit Ports - TX Buffer Ports --------------------
		gt2_txbufstatus_out         : out std_logic_vector(1 downto 0);
		------------------ Transmit Ports - TX Data Path interface -----------------
		gt2_txdata_in               : in  std_logic_vector(63 downto 0);
		---------------- Transmit Ports - TX Driver and OOB signaling --------------
		gt2_gthtxn_out              : out std_logic;
		gt2_gthtxp_out              : out std_logic;
		--------------------- Transmit Ports - TX Gearbox Ports --------------------
		gt2_txsequence_in           : in  std_logic_vector(6 downto 0);
		------------- Transmit Ports - TX Initialization and Reset Ports -----------
		gt2_txpcsreset_in           : in  std_logic;
		gt2_txresetdone_out         : out std_logic;
		----------------- Transmit Ports - TX Polarity Control Ports ---------------
		gt2_txpolarity_in           : in  std_logic;
		------------------ Transmit Ports - pattern Generator Ports ----------------
		gt2_txprbssel_in            : in  std_logic_vector(2 downto 0);

		--GT3  (X0Y39)
		--____________________________CHANNEL PORTS________________________________
		---------------------------- Channel - DRP Ports  --------------------------
		gt3_drpaddr_in              : in  std_logic_vector(8 downto 0);
		gt3_drpdi_in                : in  std_logic_vector(15 downto 0);
		gt3_drpdo_out               : out std_logic_vector(15 downto 0);
		gt3_drpen_in                : in  std_logic;
		gt3_drprdy_out              : out std_logic;
		gt3_drpwe_in                : in  std_logic;
		------------------------------- Loopback Ports -----------------------------
		gt3_loopback_in             : in  std_logic_vector(2 downto 0);
		--------------------- RX Initialization and Reset Ports --------------------
		gt3_eyescanreset_in         : in  std_logic;
		gt3_rxuserrdy_in            : in  std_logic;
		-------------------------- RX Margin Analysis Ports ------------------------
		gt3_eyescandataerror_out    : out std_logic;
		gt3_eyescantrigger_in       : in  std_logic;
		------------------- Receive Ports - Digital Monitor Ports ------------------
		gt3_dmonitorout_out         : out std_logic_vector(14 downto 0);
		------------------ Receive Ports - FPGA RX interface Ports -----------------
		gt3_rxdata_out              : out std_logic_vector(63 downto 0);
		------------------- Receive Ports - Pattern Checker Ports ------------------
		gt3_rxprbserr_out           : out std_logic;
		gt3_rxprbssel_in            : in  std_logic_vector(2 downto 0);
		------------------- Receive Ports - Pattern Checker ports ------------------
		gt3_rxprbscntreset_in       : in  std_logic;
		------------------------ Receive Ports - RX AFE Ports ----------------------
		gt3_gthrxn_in               : in  std_logic;
		------------------- Receive Ports - RX Buffer Bypass Ports -----------------
		gt3_rxbufreset_in           : in  std_logic;
		gt3_rxbufstatus_out         : out std_logic_vector(2 downto 0);
		--------------------- Receive Ports - RX Equalizer Ports -------------------
		gt3_rxmonitorout_out        : out std_logic_vector(6 downto 0);
		gt3_rxmonitorsel_in         : in  std_logic_vector(1 downto 0);
		---------------------- Receive Ports - RX Gearbox Ports --------------------
		gt3_rxdatavalid_out         : out std_logic;
		gt3_rxheader_out            : out std_logic_vector(1 downto 0);
		gt3_rxheadervalid_out       : out std_logic;
		--------------------- Receive Ports - RX Gearbox Ports  --------------------
		gt3_rxgearboxslip_in        : in  std_logic;
		------------- Receive Ports - RX Initialization and Reset Ports ------------
		gt3_gtrxreset_in            : in  std_logic;
		gt3_rxpcsreset_in           : in  std_logic;
		------------------------ Receive Ports -RX AFE Ports -----------------------
		gt3_gthrxp_in               : in  std_logic;
		-------------- Receive Ports -RX Initialization and Reset Ports ------------
		gt3_rxresetdone_out         : out std_logic;
		--------------------- TX Initialization and Reset Ports --------------------
		gt3_gttxreset_in            : in  std_logic;
		gt3_txuserrdy_in            : in  std_logic;
		-------------- Transmit Ports - 64b66b and 64b67b Gearbox Ports ------------
		gt3_txheader_in             : in  std_logic_vector(1 downto 0);
		--------------------- Transmit Ports - PCI Express Ports -------------------
		gt3_txelecidle_in           : in  std_logic;
		------------------ Transmit Ports - Pattern Generator Ports ----------------
		gt3_txprbsforceerr_in       : in  std_logic;
		---------------------- Transmit Ports - TX Buffer Ports --------------------
		gt3_txbufstatus_out         : out std_logic_vector(1 downto 0);
		------------------ Transmit Ports - TX Data Path interface -----------------
		gt3_txdata_in               : in  std_logic_vector(63 downto 0);
		---------------- Transmit Ports - TX Driver and OOB signaling --------------
		gt3_gthtxn_out              : out std_logic;
		gt3_gthtxp_out              : out std_logic;
		--------------------- Transmit Ports - TX Gearbox Ports --------------------
		gt3_txsequence_in           : in  std_logic_vector(6 downto 0);
		------------- Transmit Ports - TX Initialization and Reset Ports -----------
		gt3_txpcsreset_in           : in  std_logic;
		gt3_txresetdone_out         : out std_logic;
		----------------- Transmit Ports - TX Polarity Control Ports ---------------
		gt3_txpolarity_in           : in  std_logic;
		------------------ Transmit Ports - pattern Generator Ports ----------------
		gt3_txprbssel_in            : in  std_logic_vector(2 downto 0)
	);
end XLAUI_support;

architecture RTL of XLAUI_support is
	attribute DowngradeIPIdentifiedWarnings : string;
	attribute DowngradeIPIdentifiedWarnings of RTL : architecture is "yes";

	--**************************Component Declarations*****************************
	component XLAUI
		port(
			SYSCLK_IN                   : in  std_logic;
			SOFT_RESET_IN               : in  std_logic;
			DONT_RESET_ON_DATA_ERROR_IN : in  std_logic;
			GT0_TX_FSM_RESET_DONE_OUT   : out std_logic;
			GT0_RX_FSM_RESET_DONE_OUT   : out std_logic;
			GT0_DATA_VALID_IN           : in  std_logic;
			GT0_TX_MMCM_LOCK_IN         : in  std_logic;
			GT0_TX_MMCM_RESET_OUT       : out std_logic;
			GT0_RX_MMCM_LOCK_IN         : in  std_logic;
			GT0_RX_MMCM_RESET_OUT       : out std_logic;
			GT1_TX_FSM_RESET_DONE_OUT   : out std_logic;
			GT1_RX_FSM_RESET_DONE_OUT   : out std_logic;
			GT1_DATA_VALID_IN           : in  std_logic;
			GT1_TX_MMCM_LOCK_IN         : in  std_logic;
			GT1_TX_MMCM_RESET_OUT       : out std_logic;
			GT1_RX_MMCM_LOCK_IN         : in  std_logic;
			GT1_RX_MMCM_RESET_OUT       : out std_logic;
			GT2_TX_FSM_RESET_DONE_OUT   : out std_logic;
			GT2_RX_FSM_RESET_DONE_OUT   : out std_logic;
			GT2_DATA_VALID_IN           : in  std_logic;
			GT2_TX_MMCM_LOCK_IN         : in  std_logic;
			GT2_TX_MMCM_RESET_OUT       : out std_logic;
			GT2_RX_MMCM_LOCK_IN         : in  std_logic;
			GT2_RX_MMCM_RESET_OUT       : out std_logic;
			GT3_TX_FSM_RESET_DONE_OUT   : out std_logic;
			GT3_RX_FSM_RESET_DONE_OUT   : out std_logic;
			GT3_DATA_VALID_IN           : in  std_logic;
			GT3_TX_MMCM_LOCK_IN         : in  std_logic;
			GT3_TX_MMCM_RESET_OUT       : out std_logic;
			GT3_RX_MMCM_LOCK_IN         : in  std_logic;
			GT3_RX_MMCM_RESET_OUT       : out std_logic;

			--_________________________________________________________________________
			--GT0  (X0Y36)
			--____________________________CHANNEL PORTS________________________________
			---------------------------- Channel - DRP Ports  --------------------------
			gt0_drpaddr_in              : in  std_logic_vector(8 downto 0);
			gt0_drpclk_in               : in  std_logic;
			gt0_drpdi_in                : in  std_logic_vector(15 downto 0);
			gt0_drpdo_out               : out std_logic_vector(15 downto 0);
			gt0_drpen_in                : in  std_logic;
			gt0_drprdy_out              : out std_logic;
			gt0_drpwe_in                : in  std_logic;
			------------------------------- Loopback Ports -----------------------------
			gt0_loopback_in             : in  std_logic_vector(2 downto 0);
			--------------------- RX Initialization and Reset Ports --------------------
			gt0_eyescanreset_in         : in  std_logic;
			gt0_rxuserrdy_in            : in  std_logic;
			-------------------------- RX Margin Analysis Ports ------------------------
			gt0_eyescandataerror_out    : out std_logic;
			gt0_eyescantrigger_in       : in  std_logic;
			------------------- Receive Ports - Digital Monitor Ports ------------------
			gt0_dmonitorout_out         : out std_logic_vector(14 downto 0);
			------------------ Receive Ports - FPGA RX Interface Ports -----------------
			gt0_rxusrclk_in             : in  std_logic;
			gt0_rxusrclk2_in            : in  std_logic;
			------------------ Receive Ports - FPGA RX interface Ports -----------------
			gt0_rxdata_out              : out std_logic_vector(63 downto 0);
			------------------- Receive Ports - Pattern Checker Ports ------------------
			gt0_rxprbserr_out           : out std_logic;
			gt0_rxprbssel_in            : in  std_logic_vector(2 downto 0);
			------------------- Receive Ports - Pattern Checker ports ------------------
			gt0_rxprbscntreset_in       : in  std_logic;
			------------------------ Receive Ports - RX AFE Ports ----------------------
			gt0_gthrxn_in               : in  std_logic;
			------------------- Receive Ports - RX Buffer Bypass Ports -----------------
			gt0_rxbufreset_in           : in  std_logic;
			gt0_rxbufstatus_out         : out std_logic_vector(2 downto 0);
			--------------------- Receive Ports - RX Equalizer Ports -------------------
			gt0_rxmonitorout_out        : out std_logic_vector(6 downto 0);
			gt0_rxmonitorsel_in         : in  std_logic_vector(1 downto 0);
			--------------- Receive Ports - RX Fabric Output Control Ports -------------
			gt0_rxoutclk_out            : out std_logic;
			---------------------- Receive Ports - RX Gearbox Ports --------------------
			gt0_rxdatavalid_out         : out std_logic;
			gt0_rxheader_out            : out std_logic_vector(1 downto 0);
			gt0_rxheadervalid_out       : out std_logic;
			--------------------- Receive Ports - RX Gearbox Ports  --------------------
			gt0_rxgearboxslip_in        : in  std_logic;
			------------- Receive Ports - RX Initialization and Reset Ports ------------
			gt0_gtrxreset_in            : in  std_logic;
			gt0_rxpcsreset_in           : in  std_logic;
			------------------------ Receive Ports -RX AFE Ports -----------------------
			gt0_gthrxp_in               : in  std_logic;
			-------------- Receive Ports -RX Initialization and Reset Ports ------------
			gt0_rxresetdone_out         : out std_logic;
			--------------------- TX Initialization and Reset Ports --------------------
			gt0_gttxreset_in            : in  std_logic;
			gt0_txuserrdy_in            : in  std_logic;
			-------------- Transmit Ports - 64b66b and 64b67b Gearbox Ports ------------
			gt0_txheader_in             : in  std_logic_vector(1 downto 0);
			------------------ Transmit Ports - FPGA TX Interface Ports ----------------
			gt0_txusrclk_in             : in  std_logic;
			gt0_txusrclk2_in            : in  std_logic;
			--------------------- Transmit Ports - PCI Express Ports -------------------
			gt0_txelecidle_in           : in  std_logic;
			------------------ Transmit Ports - Pattern Generator Ports ----------------
			gt0_txprbsforceerr_in       : in  std_logic;
			---------------------- Transmit Ports - TX Buffer Ports --------------------
			gt0_txbufstatus_out         : out std_logic_vector(1 downto 0);
			------------------ Transmit Ports - TX Data Path interface -----------------
			gt0_txdata_in               : in  std_logic_vector(63 downto 0);
			---------------- Transmit Ports - TX Driver and OOB signaling --------------
			gt0_gthtxn_out              : out std_logic;
			gt0_gthtxp_out              : out std_logic;
			----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
			gt0_txoutclk_out            : out std_logic;
			gt0_txoutclkfabric_out      : out std_logic;
			gt0_txoutclkpcs_out         : out std_logic;
			--------------------- Transmit Ports - TX Gearbox Ports --------------------
			gt0_txsequence_in           : in  std_logic_vector(6 downto 0);
			------------- Transmit Ports - TX Initialization and Reset Ports -----------
			gt0_txpcsreset_in           : in  std_logic;
			gt0_txresetdone_out         : out std_logic;
			----------------- Transmit Ports - TX Polarity Control Ports ---------------
			gt0_txpolarity_in           : in  std_logic;
			------------------ Transmit Ports - pattern Generator Ports ----------------
			gt0_txprbssel_in            : in  std_logic_vector(2 downto 0);

			--GT1  (X0Y37)
			--____________________________CHANNEL PORTS________________________________
			---------------------------- Channel - DRP Ports  --------------------------
			gt1_drpaddr_in              : in  std_logic_vector(8 downto 0);
			gt1_drpclk_in               : in  std_logic;
			gt1_drpdi_in                : in  std_logic_vector(15 downto 0);
			gt1_drpdo_out               : out std_logic_vector(15 downto 0);
			gt1_drpen_in                : in  std_logic;
			gt1_drprdy_out              : out std_logic;
			gt1_drpwe_in                : in  std_logic;
			------------------------------- Loopback Ports -----------------------------
			gt1_loopback_in             : in  std_logic_vector(2 downto 0);
			--------------------- RX Initialization and Reset Ports --------------------
			gt1_eyescanreset_in         : in  std_logic;
			gt1_rxuserrdy_in            : in  std_logic;
			-------------------------- RX Margin Analysis Ports ------------------------
			gt1_eyescandataerror_out    : out std_logic;
			gt1_eyescantrigger_in       : in  std_logic;
			------------------- Receive Ports - Digital Monitor Ports ------------------
			gt1_dmonitorout_out         : out std_logic_vector(14 downto 0);
			------------------ Receive Ports - FPGA RX Interface Ports -----------------
			gt1_rxusrclk_in             : in  std_logic;
			gt1_rxusrclk2_in            : in  std_logic;
			------------------ Receive Ports - FPGA RX interface Ports -----------------
			gt1_rxdata_out              : out std_logic_vector(63 downto 0);
			------------------- Receive Ports - Pattern Checker Ports ------------------
			gt1_rxprbserr_out           : out std_logic;
			gt1_rxprbssel_in            : in  std_logic_vector(2 downto 0);
			------------------- Receive Ports - Pattern Checker ports ------------------
			gt1_rxprbscntreset_in       : in  std_logic;
			------------------------ Receive Ports - RX AFE Ports ----------------------
			gt1_gthrxn_in               : in  std_logic;
			------------------- Receive Ports - RX Buffer Bypass Ports -----------------
			gt1_rxbufreset_in           : in  std_logic;
			gt1_rxbufstatus_out         : out std_logic_vector(2 downto 0);
			--------------------- Receive Ports - RX Equalizer Ports -------------------
			gt1_rxmonitorout_out        : out std_logic_vector(6 downto 0);
			gt1_rxmonitorsel_in         : in  std_logic_vector(1 downto 0);
			--------------- Receive Ports - RX Fabric Output Control Ports -------------
			gt1_rxoutclk_out            : out std_logic;
			---------------------- Receive Ports - RX Gearbox Ports --------------------
			gt1_rxdatavalid_out         : out std_logic;
			gt1_rxheader_out            : out std_logic_vector(1 downto 0);
			gt1_rxheadervalid_out       : out std_logic;
			--------------------- Receive Ports - RX Gearbox Ports  --------------------
			gt1_rxgearboxslip_in        : in  std_logic;
			------------- Receive Ports - RX Initialization and Reset Ports ------------
			gt1_gtrxreset_in            : in  std_logic;
			gt1_rxpcsreset_in           : in  std_logic;
			------------------------ Receive Ports -RX AFE Ports -----------------------
			gt1_gthrxp_in               : in  std_logic;
			-------------- Receive Ports -RX Initialization and Reset Ports ------------
			gt1_rxresetdone_out         : out std_logic;
			--------------------- TX Initialization and Reset Ports --------------------
			gt1_gttxreset_in            : in  std_logic;
			gt1_txuserrdy_in            : in  std_logic;
			-------------- Transmit Ports - 64b66b and 64b67b Gearbox Ports ------------
			gt1_txheader_in             : in  std_logic_vector(1 downto 0);
			------------------ Transmit Ports - FPGA TX Interface Ports ----------------
			gt1_txusrclk_in             : in  std_logic;
			gt1_txusrclk2_in            : in  std_logic;
			--------------------- Transmit Ports - PCI Express Ports -------------------
			gt1_txelecidle_in           : in  std_logic;
			------------------ Transmit Ports - Pattern Generator Ports ----------------
			gt1_txprbsforceerr_in       : in  std_logic;
			---------------------- Transmit Ports - TX Buffer Ports --------------------
			gt1_txbufstatus_out         : out std_logic_vector(1 downto 0);
			------------------ Transmit Ports - TX Data Path interface -----------------
			gt1_txdata_in               : in  std_logic_vector(63 downto 0);
			---------------- Transmit Ports - TX Driver and OOB signaling --------------
			gt1_gthtxn_out              : out std_logic;
			gt1_gthtxp_out              : out std_logic;
			----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
			gt1_txoutclk_out            : out std_logic;
			gt1_txoutclkfabric_out      : out std_logic;
			gt1_txoutclkpcs_out         : out std_logic;
			--------------------- Transmit Ports - TX Gearbox Ports --------------------
			gt1_txsequence_in           : in  std_logic_vector(6 downto 0);
			------------- Transmit Ports - TX Initialization and Reset Ports -----------
			gt1_txpcsreset_in           : in  std_logic;
			gt1_txresetdone_out         : out std_logic;
			----------------- Transmit Ports - TX Polarity Control Ports ---------------
			gt1_txpolarity_in           : in  std_logic;
			------------------ Transmit Ports - pattern Generator Ports ----------------
			gt1_txprbssel_in            : in  std_logic_vector(2 downto 0);

			--GT2  (X0Y38)
			--____________________________CHANNEL PORTS________________________________
			---------------------------- Channel - DRP Ports  --------------------------
			gt2_drpaddr_in              : in  std_logic_vector(8 downto 0);
			gt2_drpclk_in               : in  std_logic;
			gt2_drpdi_in                : in  std_logic_vector(15 downto 0);
			gt2_drpdo_out               : out std_logic_vector(15 downto 0);
			gt2_drpen_in                : in  std_logic;
			gt2_drprdy_out              : out std_logic;
			gt2_drpwe_in                : in  std_logic;
			------------------------------- Loopback Ports -----------------------------
			gt2_loopback_in             : in  std_logic_vector(2 downto 0);
			--------------------- RX Initialization and Reset Ports --------------------
			gt2_eyescanreset_in         : in  std_logic;
			gt2_rxuserrdy_in            : in  std_logic;
			-------------------------- RX Margin Analysis Ports ------------------------
			gt2_eyescandataerror_out    : out std_logic;
			gt2_eyescantrigger_in       : in  std_logic;
			------------------- Receive Ports - Digital Monitor Ports ------------------
			gt2_dmonitorout_out         : out std_logic_vector(14 downto 0);
			------------------ Receive Ports - FPGA RX Interface Ports -----------------
			gt2_rxusrclk_in             : in  std_logic;
			gt2_rxusrclk2_in            : in  std_logic;
			------------------ Receive Ports - FPGA RX interface Ports -----------------
			gt2_rxdata_out              : out std_logic_vector(63 downto 0);
			------------------- Receive Ports - Pattern Checker Ports ------------------
			gt2_rxprbserr_out           : out std_logic;
			gt2_rxprbssel_in            : in  std_logic_vector(2 downto 0);
			------------------- Receive Ports - Pattern Checker ports ------------------
			gt2_rxprbscntreset_in       : in  std_logic;
			------------------------ Receive Ports - RX AFE Ports ----------------------
			gt2_gthrxn_in               : in  std_logic;
			------------------- Receive Ports - RX Buffer Bypass Ports -----------------
			gt2_rxbufreset_in           : in  std_logic;
			gt2_rxbufstatus_out         : out std_logic_vector(2 downto 0);
			--------------------- Receive Ports - RX Equalizer Ports -------------------
			gt2_rxmonitorout_out        : out std_logic_vector(6 downto 0);
			gt2_rxmonitorsel_in         : in  std_logic_vector(1 downto 0);
			--------------- Receive Ports - RX Fabric Output Control Ports -------------
			gt2_rxoutclk_out            : out std_logic;
			---------------------- Receive Ports - RX Gearbox Ports --------------------
			gt2_rxdatavalid_out         : out std_logic;
			gt2_rxheader_out            : out std_logic_vector(1 downto 0);
			gt2_rxheadervalid_out       : out std_logic;
			--------------------- Receive Ports - RX Gearbox Ports  --------------------
			gt2_rxgearboxslip_in        : in  std_logic;
			------------- Receive Ports - RX Initialization and Reset Ports ------------
			gt2_gtrxreset_in            : in  std_logic;
			gt2_rxpcsreset_in           : in  std_logic;
			------------------------ Receive Ports -RX AFE Ports -----------------------
			gt2_gthrxp_in               : in  std_logic;
			-------------- Receive Ports -RX Initialization and Reset Ports ------------
			gt2_rxresetdone_out         : out std_logic;
			--------------------- TX Initialization and Reset Ports --------------------
			gt2_gttxreset_in            : in  std_logic;
			gt2_txuserrdy_in            : in  std_logic;
			-------------- Transmit Ports - 64b66b and 64b67b Gearbox Ports ------------
			gt2_txheader_in             : in  std_logic_vector(1 downto 0);
			------------------ Transmit Ports - FPGA TX Interface Ports ----------------
			gt2_txusrclk_in             : in  std_logic;
			gt2_txusrclk2_in            : in  std_logic;
			--------------------- Transmit Ports - PCI Express Ports -------------------
			gt2_txelecidle_in           : in  std_logic;
			------------------ Transmit Ports - Pattern Generator Ports ----------------
			gt2_txprbsforceerr_in       : in  std_logic;
			---------------------- Transmit Ports - TX Buffer Ports --------------------
			gt2_txbufstatus_out         : out std_logic_vector(1 downto 0);
			------------------ Transmit Ports - TX Data Path interface -----------------
			gt2_txdata_in               : in  std_logic_vector(63 downto 0);
			---------------- Transmit Ports - TX Driver and OOB signaling --------------
			gt2_gthtxn_out              : out std_logic;
			gt2_gthtxp_out              : out std_logic;
			----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
			gt2_txoutclk_out            : out std_logic;
			gt2_txoutclkfabric_out      : out std_logic;
			gt2_txoutclkpcs_out         : out std_logic;
			--------------------- Transmit Ports - TX Gearbox Ports --------------------
			gt2_txsequence_in           : in  std_logic_vector(6 downto 0);
			------------- Transmit Ports - TX Initialization and Reset Ports -----------
			gt2_txpcsreset_in           : in  std_logic;
			gt2_txresetdone_out         : out std_logic;
			----------------- Transmit Ports - TX Polarity Control Ports ---------------
			gt2_txpolarity_in           : in  std_logic;
			------------------ Transmit Ports - pattern Generator Ports ----------------
			gt2_txprbssel_in            : in  std_logic_vector(2 downto 0);

			--GT3  (X0Y39)
			--____________________________CHANNEL PORTS________________________________
			---------------------------- Channel - DRP Ports  --------------------------
			gt3_drpaddr_in              : in  std_logic_vector(8 downto 0);
			gt3_drpclk_in               : in  std_logic;
			gt3_drpdi_in                : in  std_logic_vector(15 downto 0);
			gt3_drpdo_out               : out std_logic_vector(15 downto 0);
			gt3_drpen_in                : in  std_logic;
			gt3_drprdy_out              : out std_logic;
			gt3_drpwe_in                : in  std_logic;
			------------------------------- Loopback Ports -----------------------------
			gt3_loopback_in             : in  std_logic_vector(2 downto 0);
			--------------------- RX Initialization and Reset Ports --------------------
			gt3_eyescanreset_in         : in  std_logic;
			gt3_rxuserrdy_in            : in  std_logic;
			-------------------------- RX Margin Analysis Ports ------------------------
			gt3_eyescandataerror_out    : out std_logic;
			gt3_eyescantrigger_in       : in  std_logic;
			------------------- Receive Ports - Digital Monitor Ports ------------------
			gt3_dmonitorout_out         : out std_logic_vector(14 downto 0);
			------------------ Receive Ports - FPGA RX Interface Ports -----------------
			gt3_rxusrclk_in             : in  std_logic;
			gt3_rxusrclk2_in            : in  std_logic;
			------------------ Receive Ports - FPGA RX interface Ports -----------------
			gt3_rxdata_out              : out std_logic_vector(63 downto 0);
			------------------- Receive Ports - Pattern Checker Ports ------------------
			gt3_rxprbserr_out           : out std_logic;
			gt3_rxprbssel_in            : in  std_logic_vector(2 downto 0);
			------------------- Receive Ports - Pattern Checker ports ------------------
			gt3_rxprbscntreset_in       : in  std_logic;
			------------------------ Receive Ports - RX AFE Ports ----------------------
			gt3_gthrxn_in               : in  std_logic;
			------------------- Receive Ports - RX Buffer Bypass Ports -----------------
			gt3_rxbufreset_in           : in  std_logic;
			gt3_rxbufstatus_out         : out std_logic_vector(2 downto 0);
			--------------------- Receive Ports - RX Equalizer Ports -------------------
			gt3_rxmonitorout_out        : out std_logic_vector(6 downto 0);
			gt3_rxmonitorsel_in         : in  std_logic_vector(1 downto 0);
			--------------- Receive Ports - RX Fabric Output Control Ports -------------
			gt3_rxoutclk_out            : out std_logic;
			---------------------- Receive Ports - RX Gearbox Ports --------------------
			gt3_rxdatavalid_out         : out std_logic;
			gt3_rxheader_out            : out std_logic_vector(1 downto 0);
			gt3_rxheadervalid_out       : out std_logic;
			--------------------- Receive Ports - RX Gearbox Ports  --------------------
			gt3_rxgearboxslip_in        : in  std_logic;
			------------- Receive Ports - RX Initialization and Reset Ports ------------
			gt3_gtrxreset_in            : in  std_logic;
			gt3_rxpcsreset_in           : in  std_logic;
			------------------------ Receive Ports -RX AFE Ports -----------------------
			gt3_gthrxp_in               : in  std_logic;
			-------------- Receive Ports -RX Initialization and Reset Ports ------------
			gt3_rxresetdone_out         : out std_logic;
			--------------------- TX Initialization and Reset Ports --------------------
			gt3_gttxreset_in            : in  std_logic;
			gt3_txuserrdy_in            : in  std_logic;
			-------------- Transmit Ports - 64b66b and 64b67b Gearbox Ports ------------
			gt3_txheader_in             : in  std_logic_vector(1 downto 0);
			------------------ Transmit Ports - FPGA TX Interface Ports ----------------
			gt3_txusrclk_in             : in  std_logic;
			gt3_txusrclk2_in            : in  std_logic;
			--------------------- Transmit Ports - PCI Express Ports -------------------
			gt3_txelecidle_in           : in  std_logic;
			------------------ Transmit Ports - Pattern Generator Ports ----------------
			gt3_txprbsforceerr_in       : in  std_logic;
			---------------------- Transmit Ports - TX Buffer Ports --------------------
			gt3_txbufstatus_out         : out std_logic_vector(1 downto 0);
			------------------ Transmit Ports - TX Data Path interface -----------------
			gt3_txdata_in               : in  std_logic_vector(63 downto 0);
			---------------- Transmit Ports - TX Driver and OOB signaling --------------
			gt3_gthtxn_out              : out std_logic;
			gt3_gthtxp_out              : out std_logic;
			----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
			gt3_txoutclk_out            : out std_logic;
			gt3_txoutclkfabric_out      : out std_logic;
			gt3_txoutclkpcs_out         : out std_logic;
			--------------------- Transmit Ports - TX Gearbox Ports --------------------
			gt3_txsequence_in           : in  std_logic_vector(6 downto 0);
			------------- Transmit Ports - TX Initialization and Reset Ports -----------
			gt3_txpcsreset_in           : in  std_logic;
			gt3_txresetdone_out         : out std_logic;
			----------------- Transmit Ports - TX Polarity Control Ports ---------------
			gt3_txpolarity_in           : in  std_logic;
			------------------ Transmit Ports - pattern Generator Ports ----------------
			gt3_txprbssel_in            : in  std_logic_vector(2 downto 0);

			--____________________________COMMON PORTS________________________________
			GT0_QPLLLOCK_IN             : in  std_logic;
			GT0_QPLLREFCLKLOST_IN       : in  std_logic;
			GT0_QPLLRESET_OUT           : out std_logic;
			GT0_QPLLOUTCLK_IN           : in  std_logic;
			GT0_QPLLOUTREFCLK_IN        : in  std_logic
		);
	end component;

	component XLAUI_common_reset
		generic(
			STABLE_CLOCK_PERIOD : integer := 8 -- Period of the stable clock driving this state-machine, unit is [ns]
		);
		port(
			STABLE_CLOCK : in  std_logic; --Stable Clock, either a stable clock from the PCB
			SOFT_RESET   : in  std_logic; --User Reset, can be pulled any time
			COMMON_RESET : out std_logic --Reset QPLL
		);
	end component;

	component XLAUI_common
		generic(
			-- Simulation attributes
			WRAPPER_SIM_GTRESET_SPEEDUP : string := "FALSE" -- Set to "TRUE" to speed up sim reset 
		);
		port(
			QPLLPD_IN          : in  std_logic;
			GTREFCLK0_IN       : in  std_logic;
			QPLLLOCK_OUT       : out std_logic;
			QPLLLOCKDETCLK_IN  : in  std_logic;
			QPLLOUTCLK_OUT     : out std_logic;
			QPLLOUTREFCLK_OUT  : out std_logic;
			QPLLREFCLKLOST_OUT : out std_logic;
			QPLLRESET_IN       : in  std_logic
		);
	end component;

	--************************** Register Declarations ****************************

	--**************************** Wire Declarations ******************************

	constant STARTUP_DELAY : integer := 500; --AR43482: Transceiver needs to wait for 500 ns after configuration
	constant WAIT_CYCLES   : integer := STARTUP_DELAY / STABLE_CLOCK_PERIOD; -- Number of Clock-Cycles to wait after configuration
	constant WAIT_MAX      : integer := WAIT_CYCLES + 10; -- 500 ns plus some additional margin

	signal init_wait_count : std_logic_vector(7 downto 0) := (others => '0');
	signal init_wait_done  : std_logic                    := '0';

	signal qpllpd_i : std_logic := '0';

	--____________________________COMMON PORTS________________________________
	signal gt0_qplllock_i       : std_logic;
	signal gt0_qpllrefclklost_i : std_logic;
	signal gt0_qpllreset_i      : std_logic;
	signal gt0_qpllreset_t      : std_logic;
	signal gt0_qplloutclk_i     : std_logic;
	signal gt0_qplloutrefclk_i  : std_logic;

	--*********************************Wire Declarations**********************************
	------------------------------- Global Signals -----------------------------
	signal tied_to_ground_i : std_logic;
	signal tied_to_vcc_i    : std_logic;

	signal txoutclk_mmcm0_locked_i : std_logic;
	signal rxoutclk_mmcm0_locked_i : std_logic;
	signal txoutclk_mmcm0_reset_i  : std_logic;
	signal rxoutclk_mmcm0_reset_i  : std_logic;

	------------------------------- User Clocks ---------------------------------
	signal gt_txusrclk_i  : std_logic;
	signal gt_txusrclk2_i : std_logic;
	signal gt_rxusrclk_i  : std_logic;
	signal gt_rxusrclk2_i : std_logic;

	signal gt0_txmmcm_reset_i : std_logic;
	signal gt0_rxmmcm_reset_i : std_logic;
	signal gt1_txmmcm_reset_i : std_logic;
	signal gt1_rxmmcm_reset_i : std_logic;
	signal gt2_txmmcm_reset_i : std_logic;
	signal gt2_rxmmcm_reset_i : std_logic;
	signal gt3_txmmcm_reset_i : std_logic;
	signal gt3_rxmmcm_reset_i : std_logic;
	----------------------------- Reference Clocks ----------------------------

	attribute syn_noclockbuf : boolean;
	signal gtrefclk_i : std_logic;
	attribute syn_noclockbuf of gtrefclk_i : signal is true;

	signal commonreset_i : std_logic;
--**************************** Main Body of Code *******************************
begin
	process(SYS_CLK_I)
	begin
		if rising_edge(SYS_CLK_I) then
			-- The counter starts running when configuration has finished and 
			-- the clock is stable. When its maximum count-value has been reached,
			-- the 500 ns from Answer Record 43482 have been passed.
			if init_wait_count = WAIT_MAX then
				init_wait_done <= '1';
			else
				init_wait_count <= init_wait_count + 1;
			end if;

			if (init_wait_done = '1') then
				qpllpd_i <= SOFT_RESET_IN;
			end if;
		end if;
	end process;

	--  Static signal Assigments
	tied_to_ground_i <= '0';
	tied_to_vcc_i    <= '1';

	gt0_qpllreset_t <= commonreset_i or gt0_qpllreset_i;

	--IBUFDS_GTE2
	ibufds_instq9_clk0 : IBUFDS_GTE2
		port map(
			O     => gtrefclk_i,
			ODIV2 => open,
			CEB   => SOFT_RESET_IN,
			I     => GTREFCLK_PAD_P_IN,
			IB    => GTREFCLK_PAD_N_IN
		);

	GTREFCLK_O <= gtrefclk_i;

	common0_i : XLAUI_common
		generic map(
			WRAPPER_SIM_GTRESET_SPEEDUP => EXAMPLE_SIM_GTRESET_SPEEDUP
		)
		port map(
			QPLLPD_IN          => qpllpd_i,
			GTREFCLK0_IN       => gtrefclk_i,
			QPLLLOCK_OUT       => gt0_qplllock_i,
			QPLLLOCKDETCLK_IN  => SYS_CLK_I,
			QPLLOUTCLK_OUT     => gt0_qplloutclk_i,
			QPLLOUTREFCLK_OUT  => gt0_qplloutrefclk_i,
			QPLLREFCLKLOST_OUT => gt0_qpllrefclklost_i,
			QPLLRESET_IN       => gt0_qpllreset_t
		);

	common_reset_i : XLAUI_common_reset
		generic map(
			STABLE_CLOCK_PERIOD => STABLE_CLOCK_PERIOD -- Period of the stable clock driving this state-machine, unit is [ns]
		)
		port map(
			STABLE_CLOCK => SYS_CLK_I,  --Stable Clock, either a stable clock from the PCB
			SOFT_RESET   => SOFT_RESET_IN, --User Reset, can be pulled any time
			COMMON_RESET => commonreset_i --Reset QPLL
		);

	rxoutclk_mmcm0_reset_i <= gt0_rxmmcm_reset_i or gt1_rxmmcm_reset_i or gt2_rxmmcm_reset_i or gt3_rxmmcm_reset_i;

	gt_rxusrclk2_i          <= GT_RXUSRCLK2_IN;
	gt_rxusrclk_i           <= GT_RXUSRCLK_IN;
	rxoutclk_mmcm0_locked_i <= GT_RXUSRCLK_LOCKED_IN;
	GT_RXUSRCLK_RESET_OUT   <= rxoutclk_mmcm0_reset_i;

	txoutclk_mmcm0_reset_i <= gt0_txmmcm_reset_i or gt1_txmmcm_reset_i or gt2_txmmcm_reset_i or gt3_txmmcm_reset_i;

	gt_txusrclk2_i          <= GT_TXUSRCLK2_IN;
	gt_txusrclk_i           <= GT_TXUSRCLK_IN;
	txoutclk_mmcm0_locked_i <= GT_TXUSRCLK_LOCKED_IN;

	GT_TXUSRCLK_RESET_OUT_REGISTER_proc : process(SYS_CLK_I) is
	begin
		if rising_edge(SYS_CLK_I) then	
			GT_TXUSRCLK_RESET_OUT   <= txoutclk_mmcm0_reset_i;
		end if;
	end process GT_TXUSRCLK_RESET_OUT_REGISTER_proc;
	
	XLAUI_init_i : XLAUI
		port map(
			sysclk_in                   => SYS_CLK_I,
			soft_reset_in               => SOFT_RESET_IN,
			dont_reset_on_data_error_in => DONT_RESET_ON_DATA_ERROR_IN,
			gt0_tx_mmcm_lock_in         => txoutclk_mmcm0_locked_i,
			gt0_tx_mmcm_reset_out       => gt0_txmmcm_reset_i,
			gt0_rx_mmcm_lock_in         => rxoutclk_mmcm0_locked_i,
			gt0_rx_mmcm_reset_out       => gt0_rxmmcm_reset_i,
			gt0_tx_fsm_reset_done_out   => gt0_tx_fsm_reset_done_out,
			gt0_rx_fsm_reset_done_out   => gt0_rx_fsm_reset_done_out,
			gt0_data_valid_in           => gt0_data_valid_in,
			gt1_tx_mmcm_lock_in         => txoutclk_mmcm0_locked_i,
			gt1_tx_mmcm_reset_out       => gt1_txmmcm_reset_i,
			gt1_rx_mmcm_lock_in         => rxoutclk_mmcm0_locked_i,
			gt1_rx_mmcm_reset_out       => gt1_rxmmcm_reset_i,
			gt1_tx_fsm_reset_done_out   => gt1_tx_fsm_reset_done_out,
			gt1_rx_fsm_reset_done_out   => gt1_rx_fsm_reset_done_out,
			gt1_data_valid_in           => gt1_data_valid_in,
			gt2_tx_mmcm_lock_in         => txoutclk_mmcm0_locked_i,
			gt2_tx_mmcm_reset_out       => gt2_txmmcm_reset_i,
			gt2_rx_mmcm_lock_in         => rxoutclk_mmcm0_locked_i,
			gt2_rx_mmcm_reset_out       => gt2_rxmmcm_reset_i,
			gt2_tx_fsm_reset_done_out   => gt2_tx_fsm_reset_done_out,
			gt2_rx_fsm_reset_done_out   => gt2_rx_fsm_reset_done_out,
			gt2_data_valid_in           => gt2_data_valid_in,
			gt3_tx_mmcm_lock_in         => txoutclk_mmcm0_locked_i,
			gt3_tx_mmcm_reset_out       => gt3_txmmcm_reset_i,
			gt3_rx_mmcm_lock_in         => rxoutclk_mmcm0_locked_i,
			gt3_rx_mmcm_reset_out       => gt3_rxmmcm_reset_i,
			gt3_tx_fsm_reset_done_out   => gt3_tx_fsm_reset_done_out,
			gt3_rx_fsm_reset_done_out   => gt3_rx_fsm_reset_done_out,
			gt3_data_valid_in           => gt3_data_valid_in,

			--_____________________________________________________________________
			--_____________________________________________________________________
			--GT0  (X0Y36)

			---------------------------- Channel - DRP Ports  --------------------------
			gt0_drpaddr_in              => gt0_drpaddr_in,
			gt0_drpclk_in               => SYS_CLK_I,
			gt0_drpdi_in                => gt0_drpdi_in,
			gt0_drpdo_out               => gt0_drpdo_out,
			gt0_drpen_in                => gt0_drpen_in,
			gt0_drprdy_out              => gt0_drprdy_out,
			gt0_drpwe_in                => gt0_drpwe_in,
			------------------------------- Loopback Ports -----------------------------
			gt0_loopback_in             => gt0_loopback_in,
			--------------------- RX Initialization and Reset Ports --------------------
			gt0_eyescanreset_in         => gt0_eyescanreset_in,
			gt0_rxuserrdy_in            => gt0_rxuserrdy_in,
			-------------------------- RX Margin Analysis Ports ------------------------
			gt0_eyescandataerror_out    => gt0_eyescandataerror_out,
			gt0_eyescantrigger_in       => gt0_eyescantrigger_in,
			------------------- Receive Ports - Digital Monitor Ports ------------------
			gt0_dmonitorout_out         => gt0_dmonitorout_out,
			------------------ Receive Ports - FPGA RX Interface Ports -----------------
			gt0_rxusrclk_in             => gt_rxusrclk_i,
			gt0_rxusrclk2_in            => gt_rxusrclk2_i,
			--------------- Receive Ports - RX Fabric Output Control Ports -------------
			gt0_rxoutclk_out            => GT0_RXOUTCLK_OUT,
			------------------ Receive Ports - FPGA RX interface Ports -----------------
			gt0_rxdata_out              => gt0_rxdata_out,
			------------------- Receive Ports - Pattern Checker Ports ------------------
			gt0_rxprbserr_out           => gt0_rxprbserr_out,
			gt0_rxprbssel_in            => gt0_rxprbssel_in,
			------------------- Receive Ports - Pattern Checker ports ------------------
			gt0_rxprbscntreset_in       => gt0_rxprbscntreset_in,
			------------------------ Receive Ports - RX AFE Ports ----------------------
			gt0_gthrxn_in               => gt0_gthrxn_in,
			------------------- Receive Ports - RX Buffer Bypass Ports -----------------
			gt0_rxbufreset_in           => gt0_rxbufreset_in,
			gt0_rxbufstatus_out         => gt0_rxbufstatus_out,
			--------------------- Receive Ports - RX Equalizer Ports -------------------
			gt0_rxmonitorout_out        => gt0_rxmonitorout_out,
			gt0_rxmonitorsel_in         => gt0_rxmonitorsel_in,
			---------------------- Receive Ports - RX Gearbox Ports --------------------
			gt0_rxdatavalid_out         => gt0_rxdatavalid_out,
			gt0_rxheader_out            => gt0_rxheader_out,
			gt0_rxheadervalid_out       => gt0_rxheadervalid_out,
			--------------------- Receive Ports - RX Gearbox Ports  --------------------
			gt0_rxgearboxslip_in        => gt0_rxgearboxslip_in,
			------------- Receive Ports - RX Initialization and Reset Ports ------------
			gt0_gtrxreset_in            => gt0_gtrxreset_in,
			gt0_rxpcsreset_in           => gt0_rxpcsreset_in,
			------------------------ Receive Ports -RX AFE Ports -----------------------
			gt0_gthrxp_in               => gt0_gthrxp_in,
			-------------- Receive Ports -RX Initialization and Reset Ports ------------
			gt0_rxresetdone_out         => gt0_rxresetdone_out,
			--------------------- TX Initialization and Reset Ports --------------------
			gt0_gttxreset_in            => gt0_gttxreset_in,
			gt0_txuserrdy_in            => gt0_txuserrdy_in,
			-------------- Transmit Ports - 64b66b and 64b67b Gearbox Ports ------------
			gt0_txheader_in             => gt0_txheader_in,
			------------------ Transmit Ports - FPGA TX Interface Ports ----------------
			gt0_txusrclk_in             => gt_txusrclk_i,
			gt0_txusrclk2_in            => gt_txusrclk2_i,
			--------------------- Transmit Ports - PCI Express Ports -------------------
			gt0_txelecidle_in           => gt0_txelecidle_in,
			------------------ Transmit Ports - Pattern Generator Ports ----------------
			gt0_txprbsforceerr_in       => gt0_txprbsforceerr_in,
			---------------------- Transmit Ports - TX Buffer Ports --------------------
			gt0_txbufstatus_out         => gt0_txbufstatus_out,
			------------------ Transmit Ports - TX Data Path interface -----------------
			gt0_txdata_in               => gt0_txdata_in,
			---------------- Transmit Ports - TX Driver and OOB signaling --------------
			gt0_gthtxn_out              => gt0_gthtxn_out,
			gt0_gthtxp_out              => gt0_gthtxp_out,
			----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
			gt0_txoutclk_out            => GT0_TXOUTCLK_OUT,
			gt0_txoutclkfabric_out      => open,
			gt0_txoutclkpcs_out         => open,
			--------------------- Transmit Ports - TX Gearbox Ports --------------------
			gt0_txsequence_in           => gt0_txsequence_in,
			------------- Transmit Ports - TX Initialization and Reset Ports -----------
			gt0_txpcsreset_in           => gt0_txpcsreset_in,
			gt0_txresetdone_out         => gt0_txresetdone_out,
			----------------- Transmit Ports - TX Polarity Control Ports ---------------
			gt0_txpolarity_in           => gt0_txpolarity_in,
			------------------ Transmit Ports - pattern Generator Ports ----------------
			gt0_txprbssel_in            => gt0_txprbssel_in,

			--_____________________________________________________________________
			--_____________________________________________________________________
			--GT1  (X0Y37)

			---------------------------- Channel - DRP Ports  --------------------------
			gt1_drpaddr_in              => gt1_drpaddr_in,
			gt1_drpclk_in               => SYS_CLK_I,
			gt1_drpdi_in                => gt1_drpdi_in,
			gt1_drpdo_out               => gt1_drpdo_out,
			gt1_drpen_in                => gt1_drpen_in,
			gt1_drprdy_out              => gt1_drprdy_out,
			gt1_drpwe_in                => gt1_drpwe_in,
			------------------------------- Loopback Ports -----------------------------
			gt1_loopback_in             => gt1_loopback_in,
			--------------------- RX Initialization and Reset Ports --------------------
			gt1_eyescanreset_in         => gt1_eyescanreset_in,
			gt1_rxuserrdy_in            => gt1_rxuserrdy_in,
			-------------------------- RX Margin Analysis Ports ------------------------
			gt1_eyescandataerror_out    => gt1_eyescandataerror_out,
			gt1_eyescantrigger_in       => gt1_eyescantrigger_in,
			------------------- Receive Ports - Digital Monitor Ports ------------------
			gt1_dmonitorout_out         => gt1_dmonitorout_out,
			------------------ Receive Ports - FPGA RX Interface Ports -----------------
			gt1_rxusrclk_in             => gt_rxusrclk_i,
			gt1_rxusrclk2_in            => gt_rxusrclk2_i,
			------------------ Receive Ports - FPGA RX interface Ports -----------------
			gt1_rxdata_out              => gt1_rxdata_out,
			------------------- Receive Ports - Pattern Checker Ports ------------------
			gt1_rxprbserr_out           => gt1_rxprbserr_out,
			gt1_rxprbssel_in            => gt1_rxprbssel_in,
			------------------- Receive Ports - Pattern Checker ports ------------------
			gt1_rxprbscntreset_in       => gt1_rxprbscntreset_in,
			------------------------ Receive Ports - RX AFE Ports ----------------------
			gt1_gthrxn_in               => gt1_gthrxn_in,
			------------------- Receive Ports - RX Buffer Bypass Ports -----------------
			gt1_rxbufreset_in           => gt1_rxbufreset_in,
			gt1_rxbufstatus_out         => gt1_rxbufstatus_out,
			--------------------- Receive Ports - RX Equalizer Ports -------------------
			gt1_rxmonitorout_out        => gt1_rxmonitorout_out,
			gt1_rxmonitorsel_in         => gt1_rxmonitorsel_in,
			--------------- Receive Ports - RX Fabric Output Control Ports -------------
			gt1_rxoutclk_out            => open,
			---------------------- Receive Ports - RX Gearbox Ports --------------------
			gt1_rxdatavalid_out         => gt1_rxdatavalid_out,
			gt1_rxheader_out            => gt1_rxheader_out,
			gt1_rxheadervalid_out       => gt1_rxheadervalid_out,
			--------------------- Receive Ports - RX Gearbox Ports  --------------------
			gt1_rxgearboxslip_in        => gt1_rxgearboxslip_in,
			------------- Receive Ports - RX Initialization and Reset Ports ------------
			gt1_gtrxreset_in            => gt1_gtrxreset_in,
			gt1_rxpcsreset_in           => gt1_rxpcsreset_in,
			------------------------ Receive Ports -RX AFE Ports -----------------------
			gt1_gthrxp_in               => gt1_gthrxp_in,
			-------------- Receive Ports -RX Initialization and Reset Ports ------------
			gt1_rxresetdone_out         => gt1_rxresetdone_out,
			--------------------- TX Initialization and Reset Ports --------------------
			gt1_gttxreset_in            => gt1_gttxreset_in,
			gt1_txuserrdy_in            => gt1_txuserrdy_in,
			-------------- Transmit Ports - 64b66b and 64b67b Gearbox Ports ------------
			gt1_txheader_in             => gt1_txheader_in,
			------------------ Transmit Ports - FPGA TX Interface Ports ----------------
			gt1_txusrclk_in             => gt_txusrclk_i,
			gt1_txusrclk2_in            => gt_txusrclk2_i,
			--------------------- Transmit Ports - PCI Express Ports -------------------
			gt1_txelecidle_in           => gt1_txelecidle_in,
			------------------ Transmit Ports - Pattern Generator Ports ----------------
			gt1_txprbsforceerr_in       => gt1_txprbsforceerr_in,
			---------------------- Transmit Ports - TX Buffer Ports --------------------
			gt1_txbufstatus_out         => gt1_txbufstatus_out,
			------------------ Transmit Ports - TX Data Path interface -----------------
			gt1_txdata_in               => gt1_txdata_in,
			---------------- Transmit Ports - TX Driver and OOB signaling --------------
			gt1_gthtxn_out              => gt1_gthtxn_out,
			gt1_gthtxp_out              => gt1_gthtxp_out,
			----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
			gt1_txoutclk_out            => open,
			gt1_txoutclkfabric_out      => open,
			gt1_txoutclkpcs_out         => open,
			--------------------- Transmit Ports - TX Gearbox Ports --------------------
			gt1_txsequence_in           => gt1_txsequence_in,
			------------- Transmit Ports - TX Initialization and Reset Ports -----------
			gt1_txpcsreset_in           => gt1_txpcsreset_in,
			gt1_txresetdone_out         => gt1_txresetdone_out,
			----------------- Transmit Ports - TX Polarity Control Ports ---------------
			gt1_txpolarity_in           => gt1_txpolarity_in,
			------------------ Transmit Ports - pattern Generator Ports ----------------
			gt1_txprbssel_in            => gt1_txprbssel_in,

			--_____________________________________________________________________
			--_____________________________________________________________________
			--GT2  (X0Y38)

			---------------------------- Channel - DRP Ports  --------------------------
			gt2_drpaddr_in              => gt2_drpaddr_in,
			gt2_drpclk_in               => SYS_CLK_I,
			gt2_drpdi_in                => gt2_drpdi_in,
			gt2_drpdo_out               => gt2_drpdo_out,
			gt2_drpen_in                => gt2_drpen_in,
			gt2_drprdy_out              => gt2_drprdy_out,
			gt2_drpwe_in                => gt2_drpwe_in,
			------------------------------- Loopback Ports -----------------------------
			gt2_loopback_in             => gt2_loopback_in,
			--------------------- RX Initialization and Reset Ports --------------------
			gt2_eyescanreset_in         => gt2_eyescanreset_in,
			gt2_rxuserrdy_in            => gt2_rxuserrdy_in,
			-------------------------- RX Margin Analysis Ports ------------------------
			gt2_eyescandataerror_out    => gt2_eyescandataerror_out,
			gt2_eyescantrigger_in       => gt2_eyescantrigger_in,
			------------------- Receive Ports - Digital Monitor Ports ------------------
			gt2_dmonitorout_out         => gt2_dmonitorout_out,
			------------------ Receive Ports - FPGA RX Interface Ports -----------------
			gt2_rxusrclk_in             => gt_rxusrclk_i,
			gt2_rxusrclk2_in            => gt_rxusrclk2_i,
			------------------ Receive Ports - FPGA RX interface Ports -----------------
			gt2_rxdata_out              => gt2_rxdata_out,
			------------------- Receive Ports - Pattern Checker Ports ------------------
			gt2_rxprbserr_out           => gt2_rxprbserr_out,
			gt2_rxprbssel_in            => gt2_rxprbssel_in,
			------------------- Receive Ports - Pattern Checker ports ------------------
			gt2_rxprbscntreset_in       => gt2_rxprbscntreset_in,
			------------------------ Receive Ports - RX AFE Ports ----------------------
			gt2_gthrxn_in               => gt2_gthrxn_in,
			------------------- Receive Ports - RX Buffer Bypass Ports -----------------
			gt2_rxbufreset_in           => gt2_rxbufreset_in,
			gt2_rxbufstatus_out         => gt2_rxbufstatus_out,
			--------------------- Receive Ports - RX Equalizer Ports -------------------
			gt2_rxmonitorout_out        => gt2_rxmonitorout_out,
			gt2_rxmonitorsel_in         => gt2_rxmonitorsel_in,
			--------------- Receive Ports - RX Fabric Output Control Ports -------------
			gt2_rxoutclk_out            => open,
			---------------------- Receive Ports - RX Gearbox Ports --------------------
			gt2_rxdatavalid_out         => gt2_rxdatavalid_out,
			gt2_rxheader_out            => gt2_rxheader_out,
			gt2_rxheadervalid_out       => gt2_rxheadervalid_out,
			--------------------- Receive Ports - RX Gearbox Ports  --------------------
			gt2_rxgearboxslip_in        => gt2_rxgearboxslip_in,
			------------- Receive Ports - RX Initialization and Reset Ports ------------
			gt2_gtrxreset_in            => gt2_gtrxreset_in,
			gt2_rxpcsreset_in           => gt2_rxpcsreset_in,
			------------------------ Receive Ports -RX AFE Ports -----------------------
			gt2_gthrxp_in               => gt2_gthrxp_in,
			-------------- Receive Ports -RX Initialization and Reset Ports ------------
			gt2_rxresetdone_out         => gt2_rxresetdone_out,
			--------------------- TX Initialization and Reset Ports --------------------
			gt2_gttxreset_in            => gt2_gttxreset_in,
			gt2_txuserrdy_in            => gt2_txuserrdy_in,
			-------------- Transmit Ports - 64b66b and 64b67b Gearbox Ports ------------
			gt2_txheader_in             => gt2_txheader_in,
			------------------ Transmit Ports - FPGA TX Interface Ports ----------------
			gt2_txusrclk_in             => gt_txusrclk_i,
			gt2_txusrclk2_in            => gt_txusrclk2_i,
			--------------------- Transmit Ports - PCI Express Ports -------------------
			gt2_txelecidle_in           => gt2_txelecidle_in,
			------------------ Transmit Ports - Pattern Generator Ports ----------------
			gt2_txprbsforceerr_in       => gt2_txprbsforceerr_in,
			---------------------- Transmit Ports - TX Buffer Ports --------------------
			gt2_txbufstatus_out         => gt2_txbufstatus_out,
			------------------ Transmit Ports - TX Data Path interface -----------------
			gt2_txdata_in               => gt2_txdata_in,
			---------------- Transmit Ports - TX Driver and OOB signaling --------------
			gt2_gthtxn_out              => gt2_gthtxn_out,
			gt2_gthtxp_out              => gt2_gthtxp_out,
			----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
			gt2_txoutclk_out            => open,
			gt2_txoutclkfabric_out      => open,
			gt2_txoutclkpcs_out         => open,
			--------------------- Transmit Ports - TX Gearbox Ports --------------------
			gt2_txsequence_in           => gt2_txsequence_in,
			------------- Transmit Ports - TX Initialization and Reset Ports -----------
			gt2_txpcsreset_in           => gt2_txpcsreset_in,
			gt2_txresetdone_out         => gt2_txresetdone_out,
			----------------- Transmit Ports - TX Polarity Control Ports ---------------
			gt2_txpolarity_in           => gt2_txpolarity_in,
			------------------ Transmit Ports - pattern Generator Ports ----------------
			gt2_txprbssel_in            => gt2_txprbssel_in,

			--_____________________________________________________________________
			--_____________________________________________________________________
			--GT3  (X0Y39)

			---------------------------- Channel - DRP Ports  --------------------------
			gt3_drpaddr_in              => gt3_drpaddr_in,
			gt3_drpclk_in               => SYS_CLK_I,
			gt3_drpdi_in                => gt3_drpdi_in,
			gt3_drpdo_out               => gt3_drpdo_out,
			gt3_drpen_in                => gt3_drpen_in,
			gt3_drprdy_out              => gt3_drprdy_out,
			gt3_drpwe_in                => gt3_drpwe_in,
			------------------------------- Loopback Ports -----------------------------
			gt3_loopback_in             => gt3_loopback_in,
			--------------------- RX Initialization and Reset Ports --------------------
			gt3_eyescanreset_in         => gt3_eyescanreset_in,
			gt3_rxuserrdy_in            => gt3_rxuserrdy_in,
			-------------------------- RX Margin Analysis Ports ------------------------
			gt3_eyescandataerror_out    => gt3_eyescandataerror_out,
			gt3_eyescantrigger_in       => gt3_eyescantrigger_in,
			------------------- Receive Ports - Digital Monitor Ports ------------------
			gt3_dmonitorout_out         => gt3_dmonitorout_out,
			------------------ Receive Ports - FPGA RX Interface Ports -----------------
			gt3_rxusrclk_in             => gt_rxusrclk_i,
			gt3_rxusrclk2_in            => gt_rxusrclk2_i,
			------------------ Receive Ports - FPGA RX interface Ports -----------------
			gt3_rxdata_out              => gt3_rxdata_out,
			------------------- Receive Ports - Pattern Checker Ports ------------------
			gt3_rxprbserr_out           => gt3_rxprbserr_out,
			gt3_rxprbssel_in            => gt3_rxprbssel_in,
			------------------- Receive Ports - Pattern Checker ports ------------------
			gt3_rxprbscntreset_in       => gt3_rxprbscntreset_in,
			------------------------ Receive Ports - RX AFE Ports ----------------------
			gt3_gthrxn_in               => gt3_gthrxn_in,
			------------------- Receive Ports - RX Buffer Bypass Ports -----------------
			gt3_rxbufreset_in           => gt3_rxbufreset_in,
			gt3_rxbufstatus_out         => gt3_rxbufstatus_out,
			--------------------- Receive Ports - RX Equalizer Ports -------------------
			gt3_rxmonitorout_out        => gt3_rxmonitorout_out,
			gt3_rxmonitorsel_in         => gt3_rxmonitorsel_in,
			--------------- Receive Ports - RX Fabric Output Control Ports -------------
			gt3_rxoutclk_out            => open,
			---------------------- Receive Ports - RX Gearbox Ports --------------------
			gt3_rxdatavalid_out         => gt3_rxdatavalid_out,
			gt3_rxheader_out            => gt3_rxheader_out,
			gt3_rxheadervalid_out       => gt3_rxheadervalid_out,
			--------------------- Receive Ports - RX Gearbox Ports  --------------------
			gt3_rxgearboxslip_in        => gt3_rxgearboxslip_in,
			------------- Receive Ports - RX Initialization and Reset Ports ------------
			gt3_gtrxreset_in            => gt3_gtrxreset_in,
			gt3_rxpcsreset_in           => gt3_rxpcsreset_in,
			------------------------ Receive Ports -RX AFE Ports -----------------------
			gt3_gthrxp_in               => gt3_gthrxp_in,
			-------------- Receive Ports -RX Initialization and Reset Ports ------------
			gt3_rxresetdone_out         => gt3_rxresetdone_out,
			--------------------- TX Initialization and Reset Ports --------------------
			gt3_gttxreset_in            => gt3_gttxreset_in,
			gt3_txuserrdy_in            => gt3_txuserrdy_in,
			-------------- Transmit Ports - 64b66b and 64b67b Gearbox Ports ------------
			gt3_txheader_in             => gt3_txheader_in,
			------------------ Transmit Ports - FPGA TX Interface Ports ----------------
			gt3_txusrclk_in             => gt_txusrclk_i,
			gt3_txusrclk2_in            => gt_txusrclk2_i,
			--------------------- Transmit Ports - PCI Express Ports -------------------
			gt3_txelecidle_in           => gt3_txelecidle_in,
			------------------ Transmit Ports - Pattern Generator Ports ----------------
			gt3_txprbsforceerr_in       => gt3_txprbsforceerr_in,
			---------------------- Transmit Ports - TX Buffer Ports --------------------
			gt3_txbufstatus_out         => gt3_txbufstatus_out,
			------------------ Transmit Ports - TX Data Path interface -----------------
			gt3_txdata_in               => gt3_txdata_in,
			---------------- Transmit Ports - TX Driver and OOB signaling --------------
			gt3_gthtxn_out              => gt3_gthtxn_out,
			gt3_gthtxp_out              => gt3_gthtxp_out,
			----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
			gt3_txoutclk_out            => open,
			gt3_txoutclkfabric_out      => open,
			gt3_txoutclkpcs_out         => open,
			--------------------- Transmit Ports - TX Gearbox Ports --------------------
			gt3_txsequence_in           => gt3_txsequence_in,
			------------- Transmit Ports - TX Initialization and Reset Ports -----------
			gt3_txpcsreset_in           => gt3_txpcsreset_in,
			gt3_txresetdone_out         => gt3_txresetdone_out,
			----------------- Transmit Ports - TX Polarity Control Ports ---------------
			gt3_txpolarity_in           => gt3_txpolarity_in,
			------------------ Transmit Ports - pattern Generator Ports ----------------
			gt3_txprbssel_in            => gt3_txprbssel_in,
			gt0_qplllock_in             => gt0_qplllock_i,
			gt0_qpllrefclklost_in       => gt0_qpllrefclklost_i,
			gt0_qpllreset_out           => gt0_qpllreset_i,
			gt0_qplloutclk_in           => gt0_qplloutclk_i,
			gt0_qplloutrefclk_in        => gt0_qplloutrefclk_i
		);

end RTL;
