//------------------------------------------------------------------------------
//   ____  ____
//  /   /\/   /
// /___/  \  /    Vendor: Xilinx
// \   \   \/     Version : 3.3
//  \   \         Application : 7 Series FPGAs Transceivers Wizard 
//  /   /         Filename : gtwizard_0_init.v
// /___/   /\      
// \   \  /  \ 
//  \___\/\___\
//
//  Description : This module instantiates the modules required for
//                reset and initialisation of the Transceiver
//
// Module gtwizard_0_init
// Generated by Xilinx 7 Series FPGAs Transceivers Wizard
// 
// 
// (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES. 


`timescale 1ns / 1ps
`define DLY #1

//***********************************Entity Declaration************************
(* DowngradeIPIdentifiedWarnings="yes" *)
module gtwizard_0_init #
(
    parameter EXAMPLE_SIM_GTRESET_SPEEDUP            = "TRUE",     // Simulation setting for GT SecureIP model
    parameter EXAMPLE_SIMULATION                     =  0,         // Set to 1 for simulation
    parameter STABLE_CLOCK_PERIOD                    = 16,         //Period of the stable clock driving this state-machine, unit is [ns]
    parameter EXAMPLE_USE_CHIPSCOPE                  =  0          // Set to 1 to use Chipscope to drive resets

)
(
    //RR added these
input rx8b10b_en,
input tx8b10b_en,
    //RR added these PPM controller ports
input                 TX_PPM_EN,
input     [4:0]      TX_PPM_CTRL,
input                INV_TXOUT,

input           sysclk_in,
input           soft_reset_in,
input           dont_reset_on_data_error_in,
output          gt0_tx_fsm_reset_done_out,
output          gt0_rx_fsm_reset_done_out,
input           gt0_data_valid_in,
output          gt1_tx_fsm_reset_done_out,
output          gt1_rx_fsm_reset_done_out,
input           gt1_data_valid_in,
output          gt2_tx_fsm_reset_done_out,
output          gt2_rx_fsm_reset_done_out,
input           gt2_data_valid_in,
output          gt3_tx_fsm_reset_done_out,
output          gt3_rx_fsm_reset_done_out,
input           gt3_data_valid_in,
output          gt4_tx_fsm_reset_done_out,
output          gt4_rx_fsm_reset_done_out,
input           gt4_data_valid_in,
output          gt5_tx_fsm_reset_done_out,
output          gt5_rx_fsm_reset_done_out,
input           gt5_data_valid_in,
output          gt6_tx_fsm_reset_done_out,
output          gt6_rx_fsm_reset_done_out,
input           gt6_data_valid_in,
output          gt7_tx_fsm_reset_done_out,
output          gt7_rx_fsm_reset_done_out,
input           gt7_data_valid_in,
output          gt8_tx_fsm_reset_done_out,
output          gt8_rx_fsm_reset_done_out,
input           gt8_data_valid_in,
output          gt9_tx_fsm_reset_done_out,
output          gt9_rx_fsm_reset_done_out,
input           gt9_data_valid_in,

    //_________________________________________________________________________
    //GT0  (X1Y28)
    //____________________________CHANNEL PORTS________________________________
    //-------------------------- Channel - DRP Ports  --------------------------
    input   [8:0]   gt0_drpaddr_in,
    input           gt0_drpclk_in,
    input   [15:0]  gt0_drpdi_in,
    output  [15:0]  gt0_drpdo_out,
    input           gt0_drpen_in,
    output          gt0_drprdy_out,
    input           gt0_drpwe_in,
    //------------------- RX Initialization and Reset Ports --------------------
    input           gt0_eyescanreset_in,
    input           gt0_rxuserrdy_in,
    //------------------------ RX Margin Analysis Ports ------------------------
    output          gt0_eyescandataerror_out,
    input           gt0_eyescantrigger_in,
    //----------------- Receive Ports - Digital Monitor Ports ------------------
    output  [14:0]  gt0_dmonitorout_out,
    //---------------- Receive Ports - FPGA RX Interface Ports -----------------
    input           gt0_rxusrclk_in,
    input           gt0_rxusrclk2_in,
    //---------------- Receive Ports - FPGA RX interface Ports -----------------
    output  [31:0]  gt0_rxdata_out,
    //----------------- Receive Ports - Pattern Checker Ports ------------------
    output          gt0_rxprbserr_out,
    input   [2:0]   gt0_rxprbssel_in,
    //----------------- Receive Ports - Pattern Checker ports ------------------
    input           gt0_rxprbscntreset_in,
    //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
    output  [3:0]   gt0_rxdisperr_out,
    output  [3:0]   gt0_rxnotintable_out,
    //---------------------- Receive Ports - RX AFE Ports ----------------------
    input           gt0_gthrxn_in,
    //------------ Receive Ports - RX Byte and Word Alignment Ports ------------
    input           gt0_rxmcommaalignen_in,
    input           gt0_rxpcommaalignen_in,
    //---------------- Receive Ports - RX Channel Bonding Ports ----------------
    output          gt0_rxchanbondseq_out,
    input           gt0_rxchbonden_in,
    input   [2:0]   gt0_rxchbondlevel_in,
    input           gt0_rxchbondmaster_in,
    output  [4:0]   gt0_rxchbondo_out,
    input           gt0_rxchbondslave_in,
    //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
    output          gt0_rxchanisaligned_out,
    output          gt0_rxchanrealign_out,
    //------------------- Receive Ports - RX Equalizer Ports -------------------
    output  [6:0]   gt0_rxmonitorout_out,
    input   [1:0]   gt0_rxmonitorsel_in,
    //----------- Receive Ports - RX Initialization and Reset Ports ------------
    input           gt0_gtrxreset_in,
    //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    output  [3:0]   gt0_rxcharisk_out,
    //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
    input   [4:0]   gt0_rxchbondi_in,
    //---------------------- Receive Ports -RX AFE Ports -----------------------
    input           gt0_gthrxp_in,
    //------------ Receive Ports -RX Initialization and Reset Ports ------------
    output          gt0_rxresetdone_out,
    //------------------- TX Initialization and Reset Ports --------------------
    input           gt0_gttxreset_in,
    input           gt0_txuserrdy_in,
    //-------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    input   [3:0]   gt0_txchardispmode_in,
    input   [3:0]   gt0_txchardispval_in,
    //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
    input           gt0_txusrclk_in,
    input           gt0_txusrclk2_in,
    //---------------- Transmit Ports - Pattern Generator Ports ----------------
    input           gt0_txprbsforceerr_in,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [31:0]  gt0_txdata_in,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          gt0_gthtxn_out,
    output          gt0_gthtxp_out,
    //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    output          gt0_txoutclk_out,
    output          gt0_txoutclkfabric_out,
    output          gt0_txoutclkpcs_out,
    //----------- Transmit Ports - TX Initialization and Reset Ports -----------
    output          gt0_txresetdone_out,
    //---------------- Transmit Ports - pattern Generator Ports ----------------
    input   [2:0]   gt0_txprbssel_in,
    //--------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    input   [3:0]   gt0_txcharisk_in,

    //GT1  (X1Y29)
    //____________________________CHANNEL PORTS________________________________
    //-------------------------- Channel - DRP Ports  --------------------------
    input   [8:0]   gt1_drpaddr_in,
    input           gt1_drpclk_in,
    input   [15:0]  gt1_drpdi_in,
    output  [15:0]  gt1_drpdo_out,
    input           gt1_drpen_in,
    output          gt1_drprdy_out,
    input           gt1_drpwe_in,
    //------------------- RX Initialization and Reset Ports --------------------
    input           gt1_eyescanreset_in,
    input           gt1_rxuserrdy_in,
    //------------------------ RX Margin Analysis Ports ------------------------
    output          gt1_eyescandataerror_out,
    input           gt1_eyescantrigger_in,
    //----------------- Receive Ports - Digital Monitor Ports ------------------
    output  [14:0]  gt1_dmonitorout_out,
    //---------------- Receive Ports - FPGA RX Interface Ports -----------------
    input           gt1_rxusrclk_in,
    input           gt1_rxusrclk2_in,
    //---------------- Receive Ports - FPGA RX interface Ports -----------------
    output  [31:0]  gt1_rxdata_out,
    //----------------- Receive Ports - Pattern Checker Ports ------------------
    output          gt1_rxprbserr_out,
    input   [2:0]   gt1_rxprbssel_in,
    //----------------- Receive Ports - Pattern Checker ports ------------------
    input           gt1_rxprbscntreset_in,
    //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
    output  [3:0]   gt1_rxdisperr_out,
    output  [3:0]   gt1_rxnotintable_out,
    //---------------------- Receive Ports - RX AFE Ports ----------------------
    input           gt1_gthrxn_in,
    //------------ Receive Ports - RX Byte and Word Alignment Ports ------------
    input           gt1_rxmcommaalignen_in,
    input           gt1_rxpcommaalignen_in,
    //---------------- Receive Ports - RX Channel Bonding Ports ----------------
    output          gt1_rxchanbondseq_out,
    input           gt1_rxchbonden_in,
    input   [2:0]   gt1_rxchbondlevel_in,
    input           gt1_rxchbondmaster_in,
    output  [4:0]   gt1_rxchbondo_out,
    input           gt1_rxchbondslave_in,
    //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
    output          gt1_rxchanisaligned_out,
    output          gt1_rxchanrealign_out,
    //------------------- Receive Ports - RX Equalizer Ports -------------------
    output  [6:0]   gt1_rxmonitorout_out,
    input   [1:0]   gt1_rxmonitorsel_in,
    //----------- Receive Ports - RX Initialization and Reset Ports ------------
    input           gt1_gtrxreset_in,
    //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    output  [3:0]   gt1_rxcharisk_out,
    //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
    input   [4:0]   gt1_rxchbondi_in,
    //---------------------- Receive Ports -RX AFE Ports -----------------------
    input           gt1_gthrxp_in,
    //------------ Receive Ports -RX Initialization and Reset Ports ------------
    output          gt1_rxresetdone_out,
    //------------------- TX Initialization and Reset Ports --------------------
    input           gt1_gttxreset_in,
    input           gt1_txuserrdy_in,
    //-------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    input   [3:0]   gt1_txchardispmode_in,
    input   [3:0]   gt1_txchardispval_in,
    //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
    input           gt1_txusrclk_in,
    input           gt1_txusrclk2_in,
    //---------------- Transmit Ports - Pattern Generator Ports ----------------
    input           gt1_txprbsforceerr_in,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [31:0]  gt1_txdata_in,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          gt1_gthtxn_out,
    output          gt1_gthtxp_out,
    //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    output          gt1_txoutclk_out,
    output          gt1_txoutclkfabric_out,
    output          gt1_txoutclkpcs_out,
    //----------- Transmit Ports - TX Initialization and Reset Ports -----------
    output          gt1_txresetdone_out,
    //---------------- Transmit Ports - pattern Generator Ports ----------------
    input   [2:0]   gt1_txprbssel_in,
    //--------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    input   [3:0]   gt1_txcharisk_in,

    //GT2  (X1Y32)
    //____________________________CHANNEL PORTS________________________________
    //-------------------------- Channel - DRP Ports  --------------------------
    input   [8:0]   gt2_drpaddr_in,
    input           gt2_drpclk_in,
    input   [15:0]  gt2_drpdi_in,
    output  [15:0]  gt2_drpdo_out,
    input           gt2_drpen_in,
    output          gt2_drprdy_out,
    input           gt2_drpwe_in,
    //------------------- RX Initialization and Reset Ports --------------------
    input           gt2_eyescanreset_in,
    input           gt2_rxuserrdy_in,
    //------------------------ RX Margin Analysis Ports ------------------------
    output          gt2_eyescandataerror_out,
    input           gt2_eyescantrigger_in,
    //----------------- Receive Ports - Digital Monitor Ports ------------------
    output  [14:0]  gt2_dmonitorout_out,
    //---------------- Receive Ports - FPGA RX Interface Ports -----------------
    input           gt2_rxusrclk_in,
    input           gt2_rxusrclk2_in,
    //---------------- Receive Ports - FPGA RX interface Ports -----------------
    output  [31:0]  gt2_rxdata_out,
    //----------------- Receive Ports - Pattern Checker Ports ------------------
    output          gt2_rxprbserr_out,
    input   [2:0]   gt2_rxprbssel_in,
    //----------------- Receive Ports - Pattern Checker ports ------------------
    input           gt2_rxprbscntreset_in,
    //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
    output  [3:0]   gt2_rxdisperr_out,
    output  [3:0]   gt2_rxnotintable_out,
    //---------------------- Receive Ports - RX AFE Ports ----------------------
    input           gt2_gthrxn_in,
    //------------ Receive Ports - RX Byte and Word Alignment Ports ------------
    input           gt2_rxmcommaalignen_in,
    input           gt2_rxpcommaalignen_in,
    //---------------- Receive Ports - RX Channel Bonding Ports ----------------
    output          gt2_rxchanbondseq_out,
    input           gt2_rxchbonden_in,
    input   [2:0]   gt2_rxchbondlevel_in,
    input           gt2_rxchbondmaster_in,
    output  [4:0]   gt2_rxchbondo_out,
    input           gt2_rxchbondslave_in,
    //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
    output          gt2_rxchanisaligned_out,
    output          gt2_rxchanrealign_out,
    //------------------- Receive Ports - RX Equalizer Ports -------------------
    output  [6:0]   gt2_rxmonitorout_out,
    input   [1:0]   gt2_rxmonitorsel_in,
    //----------- Receive Ports - RX Initialization and Reset Ports ------------
    input           gt2_gtrxreset_in,
    //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    output  [3:0]   gt2_rxcharisk_out,
    //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
    input   [4:0]   gt2_rxchbondi_in,
    //---------------------- Receive Ports -RX AFE Ports -----------------------
    input           gt2_gthrxp_in,
    //------------ Receive Ports -RX Initialization and Reset Ports ------------
    output          gt2_rxresetdone_out,
    //------------------- TX Initialization and Reset Ports --------------------
    input           gt2_gttxreset_in,
    input           gt2_txuserrdy_in,
    //-------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    input   [3:0]   gt2_txchardispmode_in,
    input   [3:0]   gt2_txchardispval_in,
    //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
    input           gt2_txusrclk_in,
    input           gt2_txusrclk2_in,
    //---------------- Transmit Ports - Pattern Generator Ports ----------------
    input           gt2_txprbsforceerr_in,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [31:0]  gt2_txdata_in,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          gt2_gthtxn_out,
    output          gt2_gthtxp_out,
    //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    output          gt2_txoutclk_out,
    output          gt2_txoutclkfabric_out,
    output          gt2_txoutclkpcs_out,
    //----------- Transmit Ports - TX Initialization and Reset Ports -----------
    output          gt2_txresetdone_out,
    //---------------- Transmit Ports - pattern Generator Ports ----------------
    input   [2:0]   gt2_txprbssel_in,
    //--------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    input   [3:0]   gt2_txcharisk_in,

    //GT3  (X1Y33)
    //____________________________CHANNEL PORTS________________________________
    //-------------------------- Channel - DRP Ports  --------------------------
    input   [8:0]   gt3_drpaddr_in,
    input           gt3_drpclk_in,
    input   [15:0]  gt3_drpdi_in,
    output  [15:0]  gt3_drpdo_out,
    input           gt3_drpen_in,
    output          gt3_drprdy_out,
    input           gt3_drpwe_in,
    //------------------- RX Initialization and Reset Ports --------------------
    input           gt3_eyescanreset_in,
    input           gt3_rxuserrdy_in,
    //------------------------ RX Margin Analysis Ports ------------------------
    output          gt3_eyescandataerror_out,
    input           gt3_eyescantrigger_in,
    //----------------- Receive Ports - Digital Monitor Ports ------------------
    output  [14:0]  gt3_dmonitorout_out,
    //---------------- Receive Ports - FPGA RX Interface Ports -----------------
    input           gt3_rxusrclk_in,
    input           gt3_rxusrclk2_in,
    //---------------- Receive Ports - FPGA RX interface Ports -----------------
    output  [31:0]  gt3_rxdata_out,
    //----------------- Receive Ports - Pattern Checker Ports ------------------
    output          gt3_rxprbserr_out,
    input   [2:0]   gt3_rxprbssel_in,
    //----------------- Receive Ports - Pattern Checker ports ------------------
    input           gt3_rxprbscntreset_in,
    //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
    output  [3:0]   gt3_rxdisperr_out,
    output  [3:0]   gt3_rxnotintable_out,
    //---------------------- Receive Ports - RX AFE Ports ----------------------
    input           gt3_gthrxn_in,
    //------------ Receive Ports - RX Byte and Word Alignment Ports ------------
    input           gt3_rxmcommaalignen_in,
    input           gt3_rxpcommaalignen_in,
    //---------------- Receive Ports - RX Channel Bonding Ports ----------------
    output          gt3_rxchanbondseq_out,
    input           gt3_rxchbonden_in,
    input   [2:0]   gt3_rxchbondlevel_in,
    input           gt3_rxchbondmaster_in,
    output  [4:0]   gt3_rxchbondo_out,
    input           gt3_rxchbondslave_in,
    //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
    output          gt3_rxchanisaligned_out,
    output          gt3_rxchanrealign_out,
    //------------------- Receive Ports - RX Equalizer Ports -------------------
    output  [6:0]   gt3_rxmonitorout_out,
    input   [1:0]   gt3_rxmonitorsel_in,
    //----------- Receive Ports - RX Initialization and Reset Ports ------------
    input           gt3_gtrxreset_in,
    //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    output  [3:0]   gt3_rxcharisk_out,
    //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
    input   [4:0]   gt3_rxchbondi_in,
    //---------------------- Receive Ports -RX AFE Ports -----------------------
    input           gt3_gthrxp_in,
    //------------ Receive Ports -RX Initialization and Reset Ports ------------
    output          gt3_rxresetdone_out,
    //------------------- TX Initialization and Reset Ports --------------------
    input           gt3_gttxreset_in,
    input           gt3_txuserrdy_in,
    //-------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    input   [3:0]   gt3_txchardispmode_in,
    input   [3:0]   gt3_txchardispval_in,
    //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
    input           gt3_txusrclk_in,
    input           gt3_txusrclk2_in,
    //---------------- Transmit Ports - Pattern Generator Ports ----------------
    input           gt3_txprbsforceerr_in,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [31:0]  gt3_txdata_in,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          gt3_gthtxn_out,
    output          gt3_gthtxp_out,
    //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    output          gt3_txoutclk_out,
    output          gt3_txoutclkfabric_out,
    output          gt3_txoutclkpcs_out,
    //----------- Transmit Ports - TX Initialization and Reset Ports -----------
    output          gt3_txresetdone_out,
    //---------------- Transmit Ports - pattern Generator Ports ----------------
    input   [2:0]   gt3_txprbssel_in,
    //--------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    input   [3:0]   gt3_txcharisk_in,

    //GT4  (X1Y34)
    //____________________________CHANNEL PORTS________________________________
    //-------------------------- Channel - DRP Ports  --------------------------
    input   [8:0]   gt4_drpaddr_in,
    input           gt4_drpclk_in,
    input   [15:0]  gt4_drpdi_in,
    output  [15:0]  gt4_drpdo_out,
    input           gt4_drpen_in,
    output          gt4_drprdy_out,
    input           gt4_drpwe_in,
    //------------------- RX Initialization and Reset Ports --------------------
    input           gt4_eyescanreset_in,
    input           gt4_rxuserrdy_in,
    //------------------------ RX Margin Analysis Ports ------------------------
    output          gt4_eyescandataerror_out,
    input           gt4_eyescantrigger_in,
    //----------------- Receive Ports - Digital Monitor Ports ------------------
    output  [14:0]  gt4_dmonitorout_out,
    //---------------- Receive Ports - FPGA RX Interface Ports -----------------
    input           gt4_rxusrclk_in,
    input           gt4_rxusrclk2_in,
    //---------------- Receive Ports - FPGA RX interface Ports -----------------
    output  [31:0]  gt4_rxdata_out,
    //----------------- Receive Ports - Pattern Checker Ports ------------------
    output          gt4_rxprbserr_out,
    input   [2:0]   gt4_rxprbssel_in,
    //----------------- Receive Ports - Pattern Checker ports ------------------
    input           gt4_rxprbscntreset_in,
    //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
    output  [3:0]   gt4_rxdisperr_out,
    output  [3:0]   gt4_rxnotintable_out,
    //---------------------- Receive Ports - RX AFE Ports ----------------------
    input           gt4_gthrxn_in,
    //------------ Receive Ports - RX Byte and Word Alignment Ports ------------
    input           gt4_rxmcommaalignen_in,
    input           gt4_rxpcommaalignen_in,
    //---------------- Receive Ports - RX Channel Bonding Ports ----------------
    output          gt4_rxchanbondseq_out,
    input           gt4_rxchbonden_in,
    input   [2:0]   gt4_rxchbondlevel_in,
    input           gt4_rxchbondmaster_in,
    output  [4:0]   gt4_rxchbondo_out,
    input           gt4_rxchbondslave_in,
    //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
    output          gt4_rxchanisaligned_out,
    output          gt4_rxchanrealign_out,
    //------------------- Receive Ports - RX Equalizer Ports -------------------
    output  [6:0]   gt4_rxmonitorout_out,
    input   [1:0]   gt4_rxmonitorsel_in,
    //----------- Receive Ports - RX Initialization and Reset Ports ------------
    input           gt4_gtrxreset_in,
    //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    output  [3:0]   gt4_rxcharisk_out,
    //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
    input   [4:0]   gt4_rxchbondi_in,
    //---------------------- Receive Ports -RX AFE Ports -----------------------
    input           gt4_gthrxp_in,
    //------------ Receive Ports -RX Initialization and Reset Ports ------------
    output          gt4_rxresetdone_out,
    //------------------- TX Initialization and Reset Ports --------------------
    input           gt4_gttxreset_in,
    input           gt4_txuserrdy_in,
    //-------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    input   [3:0]   gt4_txchardispmode_in,
    input   [3:0]   gt4_txchardispval_in,
    //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
    input           gt4_txusrclk_in,
    input           gt4_txusrclk2_in,
    //---------------- Transmit Ports - Pattern Generator Ports ----------------
    input           gt4_txprbsforceerr_in,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [31:0]  gt4_txdata_in,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          gt4_gthtxn_out,
    output          gt4_gthtxp_out,
    //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    output          gt4_txoutclk_out,
    output          gt4_txoutclkfabric_out,
    output          gt4_txoutclkpcs_out,
    //----------- Transmit Ports - TX Initialization and Reset Ports -----------
    output          gt4_txresetdone_out,
    //---------------- Transmit Ports - pattern Generator Ports ----------------
    input   [2:0]   gt4_txprbssel_in,
    //--------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    input   [3:0]   gt4_txcharisk_in,

    //GT5  (X1Y35)
    //____________________________CHANNEL PORTS________________________________
    //-------------------------- Channel - DRP Ports  --------------------------
    input   [8:0]   gt5_drpaddr_in,
    input           gt5_drpclk_in,
    input   [15:0]  gt5_drpdi_in,
    output  [15:0]  gt5_drpdo_out,
    input           gt5_drpen_in,
    output          gt5_drprdy_out,
    input           gt5_drpwe_in,
    //------------------- RX Initialization and Reset Ports --------------------
    input           gt5_eyescanreset_in,
    input           gt5_rxuserrdy_in,
    //------------------------ RX Margin Analysis Ports ------------------------
    output          gt5_eyescandataerror_out,
    input           gt5_eyescantrigger_in,
    //----------------- Receive Ports - Digital Monitor Ports ------------------
    output  [14:0]  gt5_dmonitorout_out,
    //---------------- Receive Ports - FPGA RX Interface Ports -----------------
    input           gt5_rxusrclk_in,
    input           gt5_rxusrclk2_in,
    //---------------- Receive Ports - FPGA RX interface Ports -----------------
    output  [31:0]  gt5_rxdata_out,
    //----------------- Receive Ports - Pattern Checker Ports ------------------
    output          gt5_rxprbserr_out,
    input   [2:0]   gt5_rxprbssel_in,
    //----------------- Receive Ports - Pattern Checker ports ------------------
    input           gt5_rxprbscntreset_in,
    //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
    output  [3:0]   gt5_rxdisperr_out,
    output  [3:0]   gt5_rxnotintable_out,
    //---------------------- Receive Ports - RX AFE Ports ----------------------
    input           gt5_gthrxn_in,
    //------------ Receive Ports - RX Byte and Word Alignment Ports ------------
    input           gt5_rxmcommaalignen_in,
    input           gt5_rxpcommaalignen_in,
    //---------------- Receive Ports - RX Channel Bonding Ports ----------------
    output          gt5_rxchanbondseq_out,
    input           gt5_rxchbonden_in,
    input   [2:0]   gt5_rxchbondlevel_in,
    input           gt5_rxchbondmaster_in,
    output  [4:0]   gt5_rxchbondo_out,
    input           gt5_rxchbondslave_in,
    //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
    output          gt5_rxchanisaligned_out,
    output          gt5_rxchanrealign_out,
    //------------------- Receive Ports - RX Equalizer Ports -------------------
    output  [6:0]   gt5_rxmonitorout_out,
    input   [1:0]   gt5_rxmonitorsel_in,
    //----------- Receive Ports - RX Initialization and Reset Ports ------------
    input           gt5_gtrxreset_in,
    //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    output  [3:0]   gt5_rxcharisk_out,
    //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
    input   [4:0]   gt5_rxchbondi_in,
    //---------------------- Receive Ports -RX AFE Ports -----------------------
    input           gt5_gthrxp_in,
    //------------ Receive Ports -RX Initialization and Reset Ports ------------
    output          gt5_rxresetdone_out,
    //------------------- TX Initialization and Reset Ports --------------------
    input           gt5_gttxreset_in,
    input           gt5_txuserrdy_in,
    //-------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    input   [3:0]   gt5_txchardispmode_in,
    input   [3:0]   gt5_txchardispval_in,
    //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
    input           gt5_txusrclk_in,
    input           gt5_txusrclk2_in,
    //---------------- Transmit Ports - Pattern Generator Ports ----------------
    input           gt5_txprbsforceerr_in,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [31:0]  gt5_txdata_in,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          gt5_gthtxn_out,
    output          gt5_gthtxp_out,
    //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    output          gt5_txoutclk_out,
    output          gt5_txoutclkfabric_out,
    output          gt5_txoutclkpcs_out,
    //----------- Transmit Ports - TX Initialization and Reset Ports -----------
    output          gt5_txresetdone_out,
    //---------------- Transmit Ports - pattern Generator Ports ----------------
    input   [2:0]   gt5_txprbssel_in,
    //--------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    input   [3:0]   gt5_txcharisk_in,

    //GT6  (X1Y36)
    //____________________________CHANNEL PORTS________________________________
    //-------------------------- Channel - DRP Ports  --------------------------
    input   [8:0]   gt6_drpaddr_in,
    input           gt6_drpclk_in,
    input   [15:0]  gt6_drpdi_in,
    output  [15:0]  gt6_drpdo_out,
    input           gt6_drpen_in,
    output          gt6_drprdy_out,
    input           gt6_drpwe_in,
    //------------------- RX Initialization and Reset Ports --------------------
    input           gt6_eyescanreset_in,
    input           gt6_rxuserrdy_in,
    //------------------------ RX Margin Analysis Ports ------------------------
    output          gt6_eyescandataerror_out,
    input           gt6_eyescantrigger_in,
    //----------------- Receive Ports - Digital Monitor Ports ------------------
    output  [14:0]  gt6_dmonitorout_out,
    //---------------- Receive Ports - FPGA RX Interface Ports -----------------
    input           gt6_rxusrclk_in,
    input           gt6_rxusrclk2_in,
    //---------------- Receive Ports - FPGA RX interface Ports -----------------
    output  [31:0]  gt6_rxdata_out,
    //----------------- Receive Ports - Pattern Checker Ports ------------------
    output          gt6_rxprbserr_out,
    input   [2:0]   gt6_rxprbssel_in,
    //----------------- Receive Ports - Pattern Checker ports ------------------
    input           gt6_rxprbscntreset_in,
    //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
    output  [3:0]   gt6_rxdisperr_out,
    output  [3:0]   gt6_rxnotintable_out,
    //---------------------- Receive Ports - RX AFE Ports ----------------------
    input           gt6_gthrxn_in,
    //------------ Receive Ports - RX Byte and Word Alignment Ports ------------
    input           gt6_rxmcommaalignen_in,
    input           gt6_rxpcommaalignen_in,
    //---------------- Receive Ports - RX Channel Bonding Ports ----------------
    output          gt6_rxchanbondseq_out,
    input           gt6_rxchbonden_in,
    input   [2:0]   gt6_rxchbondlevel_in,
    input           gt6_rxchbondmaster_in,
    output  [4:0]   gt6_rxchbondo_out,
    input           gt6_rxchbondslave_in,
    //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
    output          gt6_rxchanisaligned_out,
    output          gt6_rxchanrealign_out,
    //------------------- Receive Ports - RX Equalizer Ports -------------------
    output  [6:0]   gt6_rxmonitorout_out,
    input   [1:0]   gt6_rxmonitorsel_in,
    //----------- Receive Ports - RX Initialization and Reset Ports ------------
    input           gt6_gtrxreset_in,
    //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    output  [3:0]   gt6_rxcharisk_out,
    //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
    input   [4:0]   gt6_rxchbondi_in,
    //---------------------- Receive Ports -RX AFE Ports -----------------------
    input           gt6_gthrxp_in,
    //------------ Receive Ports -RX Initialization and Reset Ports ------------
    output          gt6_rxresetdone_out,
    //------------------- TX Initialization and Reset Ports --------------------
    input           gt6_gttxreset_in,
    input           gt6_txuserrdy_in,
    //-------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    input   [3:0]   gt6_txchardispmode_in,
    input   [3:0]   gt6_txchardispval_in,
    //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
    input           gt6_txusrclk_in,
    input           gt6_txusrclk2_in,
    //---------------- Transmit Ports - Pattern Generator Ports ----------------
    input           gt6_txprbsforceerr_in,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [31:0]  gt6_txdata_in,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          gt6_gthtxn_out,
    output          gt6_gthtxp_out,
    //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    output          gt6_txoutclk_out,
    output          gt6_txoutclkfabric_out,
    output          gt6_txoutclkpcs_out,
    //----------- Transmit Ports - TX Initialization and Reset Ports -----------
    output          gt6_txresetdone_out,
    //---------------- Transmit Ports - pattern Generator Ports ----------------
    input   [2:0]   gt6_txprbssel_in,
    //--------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    input   [3:0]   gt6_txcharisk_in,

    //GT7  (X1Y37)
    //____________________________CHANNEL PORTS________________________________
    //-------------------------- Channel - DRP Ports  --------------------------
    input   [8:0]   gt7_drpaddr_in,
    input           gt7_drpclk_in,
    input   [15:0]  gt7_drpdi_in,
    output  [15:0]  gt7_drpdo_out,
    input           gt7_drpen_in,
    output          gt7_drprdy_out,
    input           gt7_drpwe_in,
    //------------------- RX Initialization and Reset Ports --------------------
    input           gt7_eyescanreset_in,
    input           gt7_rxuserrdy_in,
    //------------------------ RX Margin Analysis Ports ------------------------
    output          gt7_eyescandataerror_out,
    input           gt7_eyescantrigger_in,
    //----------------- Receive Ports - Digital Monitor Ports ------------------
    output  [14:0]  gt7_dmonitorout_out,
    //---------------- Receive Ports - FPGA RX Interface Ports -----------------
    input           gt7_rxusrclk_in,
    input           gt7_rxusrclk2_in,
    //---------------- Receive Ports - FPGA RX interface Ports -----------------
    output  [31:0]  gt7_rxdata_out,
    //----------------- Receive Ports - Pattern Checker Ports ------------------
    output          gt7_rxprbserr_out,
    input   [2:0]   gt7_rxprbssel_in,
    //----------------- Receive Ports - Pattern Checker ports ------------------
    input           gt7_rxprbscntreset_in,
    //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
    output  [3:0]   gt7_rxdisperr_out,
    output  [3:0]   gt7_rxnotintable_out,
    //---------------------- Receive Ports - RX AFE Ports ----------------------
    input           gt7_gthrxn_in,
    //------------ Receive Ports - RX Byte and Word Alignment Ports ------------
    input           gt7_rxmcommaalignen_in,
    input           gt7_rxpcommaalignen_in,
    //---------------- Receive Ports - RX Channel Bonding Ports ----------------
    output          gt7_rxchanbondseq_out,
    input           gt7_rxchbonden_in,
    input   [2:0]   gt7_rxchbondlevel_in,
    input           gt7_rxchbondmaster_in,
    output  [4:0]   gt7_rxchbondo_out,
    input           gt7_rxchbondslave_in,
    //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
    output          gt7_rxchanisaligned_out,
    output          gt7_rxchanrealign_out,
    //------------------- Receive Ports - RX Equalizer Ports -------------------
    output  [6:0]   gt7_rxmonitorout_out,
    input   [1:0]   gt7_rxmonitorsel_in,
    //----------- Receive Ports - RX Initialization and Reset Ports ------------
    input           gt7_gtrxreset_in,
    //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    output  [3:0]   gt7_rxcharisk_out,
    //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
    input   [4:0]   gt7_rxchbondi_in,
    //---------------------- Receive Ports -RX AFE Ports -----------------------
    input           gt7_gthrxp_in,
    //------------ Receive Ports -RX Initialization and Reset Ports ------------
    output          gt7_rxresetdone_out,
    //------------------- TX Initialization and Reset Ports --------------------
    input           gt7_gttxreset_in,
    input           gt7_txuserrdy_in,
    //-------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    input   [3:0]   gt7_txchardispmode_in,
    input   [3:0]   gt7_txchardispval_in,
    //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
    input           gt7_txusrclk_in,
    input           gt7_txusrclk2_in,
    //---------------- Transmit Ports - Pattern Generator Ports ----------------
    input           gt7_txprbsforceerr_in,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [31:0]  gt7_txdata_in,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          gt7_gthtxn_out,
    output          gt7_gthtxp_out,
    //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    output          gt7_txoutclk_out,
    output          gt7_txoutclkfabric_out,
    output          gt7_txoutclkpcs_out,
    //----------- Transmit Ports - TX Initialization and Reset Ports -----------
    output          gt7_txresetdone_out,
    //---------------- Transmit Ports - pattern Generator Ports ----------------
    input   [2:0]   gt7_txprbssel_in,
    //--------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    input   [3:0]   gt7_txcharisk_in,

    //GT8  (X1Y38)
    //____________________________CHANNEL PORTS________________________________
    //-------------------------- Channel - DRP Ports  --------------------------
    input   [8:0]   gt8_drpaddr_in,
    input           gt8_drpclk_in,
    input   [15:0]  gt8_drpdi_in,
    output  [15:0]  gt8_drpdo_out,
    input           gt8_drpen_in,
    output          gt8_drprdy_out,
    input           gt8_drpwe_in,
    //------------------- RX Initialization and Reset Ports --------------------
    input           gt8_eyescanreset_in,
    input           gt8_rxuserrdy_in,
    //------------------------ RX Margin Analysis Ports ------------------------
    output          gt8_eyescandataerror_out,
    input           gt8_eyescantrigger_in,
    //----------------- Receive Ports - Digital Monitor Ports ------------------
    output  [14:0]  gt8_dmonitorout_out,
    //---------------- Receive Ports - FPGA RX Interface Ports -----------------
    input           gt8_rxusrclk_in,
    input           gt8_rxusrclk2_in,
    //---------------- Receive Ports - FPGA RX interface Ports -----------------
    output  [31:0]  gt8_rxdata_out,
    //----------------- Receive Ports - Pattern Checker Ports ------------------
    output          gt8_rxprbserr_out,
    input   [2:0]   gt8_rxprbssel_in,
    //----------------- Receive Ports - Pattern Checker ports ------------------
    input           gt8_rxprbscntreset_in,
    //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
    output  [3:0]   gt8_rxdisperr_out,
    output  [3:0]   gt8_rxnotintable_out,
    //---------------------- Receive Ports - RX AFE Ports ----------------------
    input           gt8_gthrxn_in,
    //------------ Receive Ports - RX Byte and Word Alignment Ports ------------
    input           gt8_rxmcommaalignen_in,
    input           gt8_rxpcommaalignen_in,
    //---------------- Receive Ports - RX Channel Bonding Ports ----------------
    output          gt8_rxchanbondseq_out,
    input           gt8_rxchbonden_in,
    input   [2:0]   gt8_rxchbondlevel_in,
    input           gt8_rxchbondmaster_in,
    output  [4:0]   gt8_rxchbondo_out,
    input           gt8_rxchbondslave_in,
    //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
    output          gt8_rxchanisaligned_out,
    output          gt8_rxchanrealign_out,
    //------------------- Receive Ports - RX Equalizer Ports -------------------
    output  [6:0]   gt8_rxmonitorout_out,
    input   [1:0]   gt8_rxmonitorsel_in,
    //----------- Receive Ports - RX Initialization and Reset Ports ------------
    input           gt8_gtrxreset_in,
    //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    output  [3:0]   gt8_rxcharisk_out,
    //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
    input   [4:0]   gt8_rxchbondi_in,
    //---------------------- Receive Ports -RX AFE Ports -----------------------
    input           gt8_gthrxp_in,
    //------------ Receive Ports -RX Initialization and Reset Ports ------------
    output          gt8_rxresetdone_out,
    //------------------- TX Initialization and Reset Ports --------------------
    input           gt8_gttxreset_in,
    input           gt8_txuserrdy_in,
    //-------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    input   [3:0]   gt8_txchardispmode_in,
    input   [3:0]   gt8_txchardispval_in,
    //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
    input           gt8_txusrclk_in,
    input           gt8_txusrclk2_in,
    //---------------- Transmit Ports - Pattern Generator Ports ----------------
    input           gt8_txprbsforceerr_in,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [31:0]  gt8_txdata_in,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          gt8_gthtxn_out,
    output          gt8_gthtxp_out,
    //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    output          gt8_txoutclk_out,
    output          gt8_txoutclkfabric_out,
    output          gt8_txoutclkpcs_out,
    //----------- Transmit Ports - TX Initialization and Reset Ports -----------
    output          gt8_txresetdone_out,
    //---------------- Transmit Ports - pattern Generator Ports ----------------
    input   [2:0]   gt8_txprbssel_in,
    //--------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    input   [3:0]   gt8_txcharisk_in,

    //GT9  (X1Y39)
    //____________________________CHANNEL PORTS________________________________
    //-------------------------- Channel - DRP Ports  --------------------------
    input   [8:0]   gt9_drpaddr_in,
    input           gt9_drpclk_in,
    input   [15:0]  gt9_drpdi_in,
    output  [15:0]  gt9_drpdo_out,
    input           gt9_drpen_in,
    output          gt9_drprdy_out,
    input           gt9_drpwe_in,
    //------------------- RX Initialization and Reset Ports --------------------
    input           gt9_eyescanreset_in,
    input           gt9_rxuserrdy_in,
    //------------------------ RX Margin Analysis Ports ------------------------
    output          gt9_eyescandataerror_out,
    input           gt9_eyescantrigger_in,
    //----------------- Receive Ports - Digital Monitor Ports ------------------
    output  [14:0]  gt9_dmonitorout_out,
    //---------------- Receive Ports - FPGA RX Interface Ports -----------------
    input           gt9_rxusrclk_in,
    input           gt9_rxusrclk2_in,
    //---------------- Receive Ports - FPGA RX interface Ports -----------------
    output  [31:0]  gt9_rxdata_out,
    //----------------- Receive Ports - Pattern Checker Ports ------------------
    output          gt9_rxprbserr_out,
    input   [2:0]   gt9_rxprbssel_in,
    //----------------- Receive Ports - Pattern Checker ports ------------------
    input           gt9_rxprbscntreset_in,
    //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
    output  [3:0]   gt9_rxdisperr_out,
    output  [3:0]   gt9_rxnotintable_out,
    //---------------------- Receive Ports - RX AFE Ports ----------------------
    input           gt9_gthrxn_in,
    //------------ Receive Ports - RX Byte and Word Alignment Ports ------------
    input           gt9_rxmcommaalignen_in,
    input           gt9_rxpcommaalignen_in,
    //---------------- Receive Ports - RX Channel Bonding Ports ----------------
    output          gt9_rxchanbondseq_out,
    input           gt9_rxchbonden_in,
    input   [2:0]   gt9_rxchbondlevel_in,
    input           gt9_rxchbondmaster_in,
    output  [4:0]   gt9_rxchbondo_out,
    input           gt9_rxchbondslave_in,
    //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
    output          gt9_rxchanisaligned_out,
    output          gt9_rxchanrealign_out,
    //------------------- Receive Ports - RX Equalizer Ports -------------------
    output  [6:0]   gt9_rxmonitorout_out,
    input   [1:0]   gt9_rxmonitorsel_in,
    //----------- Receive Ports - RX Initialization and Reset Ports ------------
    input           gt9_gtrxreset_in,
    //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    output  [3:0]   gt9_rxcharisk_out,
    //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
    input   [4:0]   gt9_rxchbondi_in,
    //---------------------- Receive Ports -RX AFE Ports -----------------------
    input           gt9_gthrxp_in,
    //------------ Receive Ports -RX Initialization and Reset Ports ------------
    output          gt9_rxresetdone_out,
    //------------------- TX Initialization and Reset Ports --------------------
    input           gt9_gttxreset_in,
    input           gt9_txuserrdy_in,
    //-------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    input   [3:0]   gt9_txchardispmode_in,
    input   [3:0]   gt9_txchardispval_in,
    //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
    input           gt9_txusrclk_in,
    input           gt9_txusrclk2_in,
    //---------------- Transmit Ports - Pattern Generator Ports ----------------
    input           gt9_txprbsforceerr_in,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [31:0]  gt9_txdata_in,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          gt9_gthtxn_out,
    output          gt9_gthtxp_out,
    //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    output          gt9_txoutclk_out,
    output          gt9_txoutclkfabric_out,
    output          gt9_txoutclkpcs_out,
    //----------- Transmit Ports - TX Initialization and Reset Ports -----------
    output          gt9_txresetdone_out,
    //---------------- Transmit Ports - pattern Generator Ports ----------------
    input   [2:0]   gt9_txprbssel_in,
    //--------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    input   [3:0]   gt9_txcharisk_in,


    //____________________________COMMON PORTS________________________________
    input      gt0_qplllock_in,
    input      gt0_qpllrefclklost_in,
    output     gt0_qpllreset_out,
    input      gt0_qplloutclk_in,
    input      gt0_qplloutrefclk_in,
    input      gt1_qplllock_in,
    input      gt1_qpllrefclklost_in,
    output     gt1_qpllreset_out,
    input      gt1_qplloutclk_in,
    input      gt1_qplloutrefclk_in,
    input      gt2_qplllock_in,
    input      gt2_qpllrefclklost_in,
    output     gt2_qpllreset_out,
    input      gt2_qplloutclk_in,
    input      gt2_qplloutrefclk_in

);



//***********************************Parameter Declarations********************


    //Typical CDRLOCK Time is 50,000UI, as per DS183
    localparam RX_CDRLOCK_TIME      = (EXAMPLE_SIMULATION == 1) ? 1000 : 50000/10;

       
    integer   WAIT_TIME_CDRLOCK    = RX_CDRLOCK_TIME / STABLE_CLOCK_PERIOD;      

//-------------------------- GT Wrapper Wires ------------------------------
    wire           gt0_rxpmaresetdone_i;
    wire           gt0_txpmaresetdone_i;
    wire           gt0_txresetdone_i;
    wire           gt0_rxresetdone_i;
    wire           gt0_gttxreset_i;
    wire           gt0_gttxreset_t;
    wire           gt0_gtrxreset_i;
    wire           gt0_gtrxreset_t;
    wire           gt0_txuserrdy_i;
    wire           gt0_txuserrdy_t;
    wire           gt0_rxuserrdy_i;
    wire           gt0_rxuserrdy_t;

    wire           gt0_rxdfeagchold_i;
    wire           gt0_rxdfelfhold_i;
    wire           gt0_rxlpmlfhold_i;
    wire           gt0_rxlpmhfhold_i;


    wire           gt1_rxpmaresetdone_i;
    wire           gt1_txpmaresetdone_i;
    wire           gt1_txresetdone_i;
    wire           gt1_rxresetdone_i;
    wire           gt1_gttxreset_i;
    wire           gt1_gttxreset_t;
    wire           gt1_gtrxreset_i;
    wire           gt1_gtrxreset_t;
    wire           gt1_txuserrdy_i;
    wire           gt1_txuserrdy_t;
    wire           gt1_rxuserrdy_i;
    wire           gt1_rxuserrdy_t;

    wire           gt1_rxdfeagchold_i;
    wire           gt1_rxdfelfhold_i;
    wire           gt1_rxlpmlfhold_i;
    wire           gt1_rxlpmhfhold_i;


    wire           gt2_rxpmaresetdone_i;
    wire           gt2_txpmaresetdone_i;
    wire           gt2_txresetdone_i;
    wire           gt2_rxresetdone_i;
    wire           gt2_gttxreset_i;
    wire           gt2_gttxreset_t;
    wire           gt2_gtrxreset_i;
    wire           gt2_gtrxreset_t;
    wire           gt2_txuserrdy_i;
    wire           gt2_txuserrdy_t;
    wire           gt2_rxuserrdy_i;
    wire           gt2_rxuserrdy_t;

    wire           gt2_rxdfeagchold_i;
    wire           gt2_rxdfelfhold_i;
    wire           gt2_rxlpmlfhold_i;
    wire           gt2_rxlpmhfhold_i;


    wire           gt3_rxpmaresetdone_i;
    wire           gt3_txpmaresetdone_i;
    wire           gt3_txresetdone_i;
    wire           gt3_rxresetdone_i;
    wire           gt3_gttxreset_i;
    wire           gt3_gttxreset_t;
    wire           gt3_gtrxreset_i;
    wire           gt3_gtrxreset_t;
    wire           gt3_txuserrdy_i;
    wire           gt3_txuserrdy_t;
    wire           gt3_rxuserrdy_i;
    wire           gt3_rxuserrdy_t;

    wire           gt3_rxdfeagchold_i;
    wire           gt3_rxdfelfhold_i;
    wire           gt3_rxlpmlfhold_i;
    wire           gt3_rxlpmhfhold_i;


    wire           gt4_rxpmaresetdone_i;
    wire           gt4_txpmaresetdone_i;
    wire           gt4_txresetdone_i;
    wire           gt4_rxresetdone_i;
    wire           gt4_gttxreset_i;
    wire           gt4_gttxreset_t;
    wire           gt4_gtrxreset_i;
    wire           gt4_gtrxreset_t;
    wire           gt4_txuserrdy_i;
    wire           gt4_txuserrdy_t;
    wire           gt4_rxuserrdy_i;
    wire           gt4_rxuserrdy_t;

    wire           gt4_rxdfeagchold_i;
    wire           gt4_rxdfelfhold_i;
    wire           gt4_rxlpmlfhold_i;
    wire           gt4_rxlpmhfhold_i;


    wire           gt5_rxpmaresetdone_i;
    wire           gt5_txpmaresetdone_i;
    wire           gt5_txresetdone_i;
    wire           gt5_rxresetdone_i;
    wire           gt5_gttxreset_i;
    wire           gt5_gttxreset_t;
    wire           gt5_gtrxreset_i;
    wire           gt5_gtrxreset_t;
    wire           gt5_txuserrdy_i;
    wire           gt5_txuserrdy_t;
    wire           gt5_rxuserrdy_i;
    wire           gt5_rxuserrdy_t;

    wire           gt5_rxdfeagchold_i;
    wire           gt5_rxdfelfhold_i;
    wire           gt5_rxlpmlfhold_i;
    wire           gt5_rxlpmhfhold_i;


    wire           gt6_rxpmaresetdone_i;
    wire           gt6_txpmaresetdone_i;
    wire           gt6_txresetdone_i;
    wire           gt6_rxresetdone_i;
    wire           gt6_gttxreset_i;
    wire           gt6_gttxreset_t;
    wire           gt6_gtrxreset_i;
    wire           gt6_gtrxreset_t;
    wire           gt6_txuserrdy_i;
    wire           gt6_txuserrdy_t;
    wire           gt6_rxuserrdy_i;
    wire           gt6_rxuserrdy_t;

    wire           gt6_rxdfeagchold_i;
    wire           gt6_rxdfelfhold_i;
    wire           gt6_rxlpmlfhold_i;
    wire           gt6_rxlpmhfhold_i;


    wire           gt7_rxpmaresetdone_i;
    wire           gt7_txpmaresetdone_i;
    wire           gt7_txresetdone_i;
    wire           gt7_rxresetdone_i;
    wire           gt7_gttxreset_i;
    wire           gt7_gttxreset_t;
    wire           gt7_gtrxreset_i;
    wire           gt7_gtrxreset_t;
    wire           gt7_txuserrdy_i;
    wire           gt7_txuserrdy_t;
    wire           gt7_rxuserrdy_i;
    wire           gt7_rxuserrdy_t;

    wire           gt7_rxdfeagchold_i;
    wire           gt7_rxdfelfhold_i;
    wire           gt7_rxlpmlfhold_i;
    wire           gt7_rxlpmhfhold_i;


    wire           gt8_rxpmaresetdone_i;
    wire           gt8_txpmaresetdone_i;
    wire           gt8_txresetdone_i;
    wire           gt8_rxresetdone_i;
    wire           gt8_gttxreset_i;
    wire           gt8_gttxreset_t;
    wire           gt8_gtrxreset_i;
    wire           gt8_gtrxreset_t;
    wire           gt8_txuserrdy_i;
    wire           gt8_txuserrdy_t;
    wire           gt8_rxuserrdy_i;
    wire           gt8_rxuserrdy_t;

    wire           gt8_rxdfeagchold_i;
    wire           gt8_rxdfelfhold_i;
    wire           gt8_rxlpmlfhold_i;
    wire           gt8_rxlpmhfhold_i;


    wire           gt9_rxpmaresetdone_i;
    wire           gt9_txpmaresetdone_i;
    wire           gt9_txresetdone_i;
    wire           gt9_rxresetdone_i;
    wire           gt9_gttxreset_i;
    wire           gt9_gttxreset_t;
    wire           gt9_gtrxreset_i;
    wire           gt9_gtrxreset_t;
    wire           gt9_txuserrdy_i;
    wire           gt9_txuserrdy_t;
    wire           gt9_rxuserrdy_i;
    wire           gt9_rxuserrdy_t;

    wire           gt9_rxdfeagchold_i;
    wire           gt9_rxdfelfhold_i;
    wire           gt9_rxlpmlfhold_i;
    wire           gt9_rxlpmhfhold_i;



    wire           gt0_qpllreset_i;
    wire           gt0_qpllreset_t;
    wire           gt0_qpllrefclklost_i;
    wire           gt0_qplllock_i;
    wire           gt1_qpllreset_i;
    wire           gt1_qpllreset_t;
    wire           gt1_qpllrefclklost_i;
    wire           gt1_qplllock_i;
    wire           gt2_qpllreset_i;
    wire           gt2_qpllreset_t;
    wire           gt2_qpllrefclklost_i;
    wire           gt2_qplllock_i;


//------------------------------- Global Signals -----------------------------
    wire          tied_to_ground_i;
    wire          tied_to_vcc_i;

    wire           gt0_txoutclk_i;
    wire           gt0_rxoutclk_i;
    wire           gt0_rxoutclk_i2;
    wire           gt0_txoutclk_i2;
    wire           gt0_recclk_stable_i;
    reg            gt0_rx_cdrlocked;
    integer  gt0_rx_cdrlock_counter= 0;

    wire           gt1_txoutclk_i;
    wire           gt1_rxoutclk_i;
    wire           gt1_rxoutclk_i2;
    wire           gt1_txoutclk_i2;
    wire           gt1_recclk_stable_i;
    reg            gt1_rx_cdrlocked;
    integer  gt1_rx_cdrlock_counter= 0;

    wire           gt2_txoutclk_i;
    wire           gt2_rxoutclk_i;
    wire           gt2_rxoutclk_i2;
    wire           gt2_txoutclk_i2;
    wire           gt2_recclk_stable_i;
    reg            gt2_rx_cdrlocked;
    integer  gt2_rx_cdrlock_counter= 0;

    wire           gt3_txoutclk_i;
    wire           gt3_rxoutclk_i;
    wire           gt3_rxoutclk_i2;
    wire           gt3_txoutclk_i2;
    wire           gt3_recclk_stable_i;
    reg            gt3_rx_cdrlocked;
    integer  gt3_rx_cdrlock_counter= 0;

    wire           gt4_txoutclk_i;
    wire           gt4_rxoutclk_i;
    wire           gt4_rxoutclk_i2;
    wire           gt4_txoutclk_i2;
    wire           gt4_recclk_stable_i;
    reg            gt4_rx_cdrlocked;
    integer  gt4_rx_cdrlock_counter= 0;

    wire           gt5_txoutclk_i;
    wire           gt5_rxoutclk_i;
    wire           gt5_rxoutclk_i2;
    wire           gt5_txoutclk_i2;
    wire           gt5_recclk_stable_i;
    reg            gt5_rx_cdrlocked;
    integer  gt5_rx_cdrlock_counter= 0;

    wire           gt6_txoutclk_i;
    wire           gt6_rxoutclk_i;
    wire           gt6_rxoutclk_i2;
    wire           gt6_txoutclk_i2;
    wire           gt6_recclk_stable_i;
    reg            gt6_rx_cdrlocked;
    integer  gt6_rx_cdrlock_counter= 0;

    wire           gt7_txoutclk_i;
    wire           gt7_rxoutclk_i;
    wire           gt7_rxoutclk_i2;
    wire           gt7_txoutclk_i2;
    wire           gt7_recclk_stable_i;
    reg            gt7_rx_cdrlocked;
    integer  gt7_rx_cdrlock_counter= 0;

    wire           gt8_txoutclk_i;
    wire           gt8_rxoutclk_i;
    wire           gt8_rxoutclk_i2;
    wire           gt8_txoutclk_i2;
    wire           gt8_recclk_stable_i;
    reg            gt8_rx_cdrlocked;
    integer  gt8_rx_cdrlock_counter= 0;

    wire           gt9_txoutclk_i;
    wire           gt9_rxoutclk_i;
    wire           gt9_rxoutclk_i2;
    wire           gt9_txoutclk_i2;
    wire           gt9_recclk_stable_i;
    reg            gt9_rx_cdrlocked;
    integer  gt9_rx_cdrlock_counter= 0;







reg              rx_cdrlocked;


 


//**************************** Main Body of Code *******************************
    //  Static signal Assigments
assign  tied_to_ground_i                     =  1'b0;
assign  tied_to_vcc_i                        =  1'b1;

//    ----------------------------- The GT Wrapper -----------------------------
    
    // Use the instantiation template in the example directory to add the GT wrapper to your design.
    // In this example, the wrapper is wired up for basic operation with a frame generator and frame 
    // checker. The GTs will reset, then attempt to align and transmit data. If channel bonding is 
    // enabled, bonding should occur after alignment.


    gtwizard_0_multi_gt #
    (
        .EXAMPLE_SIMULATION             (EXAMPLE_SIMULATION),
        .WRAPPER_SIM_GTRESET_SPEEDUP    (EXAMPLE_SIM_GTRESET_SPEEDUP)
    )
    gtwizard_0_i
    (
        //RR added these
        .rx8b10b_en(rx8b10b_en),
        .tx8b10b_en(tx8b10b_en),
 		.TX_PPM_EN								(TX_PPM_EN),
        .TX_PPM_CTRL                            (TX_PPM_CTRL),
        .INV_TXOUT                              (INV_TXOUT),
        
         .gt0_rxpmaresetdone_out         (gt0_rxpmaresetdone_i),
        .gt0_txpmaresetdone_out         (gt0_txpmaresetdone_i),
 
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GT0  (X1Y28)

        //-------------------------- Channel - DRP Ports  --------------------------
        .gt0_drpaddr_in                 (gt0_drpaddr_in), // input wire [8:0] gt0_drpaddr_in
        .gt0_drpclk_in                  (gt0_drpclk_in), // input wire gt0_drpclk_in
        .gt0_drpdi_in                   (gt0_drpdi_in), // input wire [15:0] gt0_drpdi_in
        .gt0_drpdo_out                  (gt0_drpdo_out), // output wire [15:0] gt0_drpdo_out
        .gt0_drpen_in                   (gt0_drpen_in), // input wire gt0_drpen_in
        .gt0_drprdy_out                 (gt0_drprdy_out), // output wire gt0_drprdy_out
        .gt0_drpwe_in                   (gt0_drpwe_in), // input wire gt0_drpwe_in
        //------------------- RX Initialization and Reset Ports --------------------
        .gt0_eyescanreset_in            (gt0_eyescanreset_in), // input wire gt0_eyescanreset_in
        .gt0_rxuserrdy_in               (gt0_rxuserrdy_i), // input wire gt0_rxuserrdy_i
        //------------------------ RX Margin Analysis Ports ------------------------
        .gt0_eyescandataerror_out       (gt0_eyescandataerror_out), // output wire gt0_eyescandataerror_out
        .gt0_eyescantrigger_in          (gt0_eyescantrigger_in), // input wire gt0_eyescantrigger_in
        //----------------- Receive Ports - Digital Monitor Ports ------------------
        .gt0_dmonitorout_out            (gt0_dmonitorout_out), // output wire [14:0] gt0_dmonitorout_out
        //---------------- Receive Ports - FPGA RX Interface Ports -----------------
        .gt0_rxusrclk_in                (gt0_rxusrclk_in), // input wire gt0_rxusrclk_in
        .gt0_rxusrclk2_in               (gt0_rxusrclk2_in), // input wire gt0_rxusrclk2_in
        //---------------- Receive Ports - FPGA RX interface Ports -----------------
        .gt0_rxdata_out                 (gt0_rxdata_out), // output wire [31:0] gt0_rxdata_out
        //----------------- Receive Ports - Pattern Checker Ports ------------------
        .gt0_rxprbserr_out              (gt0_rxprbserr_out), // output wire gt0_rxprbserr_out
        .gt0_rxprbssel_in               (gt0_rxprbssel_in), // input wire [2:0] gt0_rxprbssel_in
        //----------------- Receive Ports - Pattern Checker ports ------------------
        .gt0_rxprbscntreset_in          (gt0_rxprbscntreset_in), // input wire gt0_rxprbscntreset_in
        //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
        .gt0_rxdisperr_out              (gt0_rxdisperr_out), // output wire [3:0] gt0_rxdisperr_out
        .gt0_rxnotintable_out           (gt0_rxnotintable_out), // output wire [3:0] gt0_rxnotintable_out
        //---------------------- Receive Ports - RX AFE Ports ----------------------
        .gt0_gthrxn_in                  (gt0_gthrxn_in), // input wire gt0_gthrxn_in
        //------------ Receive Ports - RX Byte and Word Alignment Ports ------------
        .gt0_rxmcommaalignen_in         (gt0_rxmcommaalignen_in), // input wire gt0_rxmcommaalignen_in
        .gt0_rxpcommaalignen_in         (gt0_rxpcommaalignen_in), // input wire gt0_rxpcommaalignen_in
        //---------------- Receive Ports - RX Channel Bonding Ports ----------------
        .gt0_rxchanbondseq_out          (gt0_rxchanbondseq_out), // output wire gt0_rxchanbondseq_out
        .gt0_rxchbonden_in              (gt0_rxchbonden_in), // input wire gt0_rxchbonden_in
        .gt0_rxchbondlevel_in           (gt0_rxchbondlevel_in), // input wire [2:0] gt0_rxchbondlevel_in
        .gt0_rxchbondmaster_in          (gt0_rxchbondmaster_in), // input wire gt0_rxchbondmaster_in
        .gt0_rxchbondo_out              (gt0_rxchbondo_out), // output wire [4:0] gt0_rxchbondo_out
        .gt0_rxchbondslave_in           (gt0_rxchbondslave_in), // input wire gt0_rxchbondslave_in
        //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
        .gt0_rxchanisaligned_out        (gt0_rxchanisaligned_out), // output wire gt0_rxchanisaligned_out
        .gt0_rxchanrealign_out          (gt0_rxchanrealign_out), // output wire gt0_rxchanrealign_out
        //------------------- Receive Ports - RX Equalizer Ports -------------------
        .gt0_rxdfeagchold_in            (gt0_rxdfeagchold_i), // input wire gt0_rxdfeagchold_i
        .gt0_rxdfelfhold_in             (gt0_rxdfelfhold_i), // input wire gt0_rxdfelfhold_i
        .gt0_rxmonitorout_out           (gt0_rxmonitorout_out), // output wire [6:0] gt0_rxmonitorout_out
        .gt0_rxmonitorsel_in            (gt0_rxmonitorsel_in), // input wire [1:0] gt0_rxmonitorsel_in
        //------------- Receive Ports - RX Fabric Output Control Ports -------------
        .gt0_rxoutclk_out               (gt0_rxoutclk_i), // output wire gt0_rxoutclk_i
        //----------- Receive Ports - RX Initialization and Reset Ports ------------
        .gt0_gtrxreset_in               (gt0_gtrxreset_i), // input wire gt0_gtrxreset_i
        //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        .gt0_rxcharisk_out              (gt0_rxcharisk_out), // output wire [3:0] gt0_rxcharisk_out
        //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
        .gt0_rxchbondi_in               (gt0_rxchbondi_in), // input wire [4:0] gt0_rxchbondi_in
        //---------------------- Receive Ports -RX AFE Ports -----------------------
        .gt0_gthrxp_in                  (gt0_gthrxp_in), // input wire gt0_gthrxp_in
        //------------ Receive Ports -RX Initialization and Reset Ports ------------
        .gt0_rxresetdone_out            (gt0_rxresetdone_i), // output wire gt0_rxresetdone_i
        //------------------- TX Initialization and Reset Ports --------------------
        .gt0_gttxreset_in               (gt0_gttxreset_i), // input wire gt0_gttxreset_i
        .gt0_txuserrdy_in               (gt0_txuserrdy_i), // input wire gt0_txuserrdy_i
        //-------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        .gt0_txchardispmode_in          (gt0_txchardispmode_in), // input wire [3:0] gt0_txchardispmode_in
        .gt0_txchardispval_in           (gt0_txchardispval_in), // input wire [3:0] gt0_txchardispval_in
        //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
        .gt0_txusrclk_in                (gt0_txusrclk_in), // input wire gt0_txusrclk_in
        .gt0_txusrclk2_in               (gt0_txusrclk2_in), // input wire gt0_txusrclk2_in
        //---------------- Transmit Ports - Pattern Generator Ports ----------------
        .gt0_txprbsforceerr_in          (gt0_txprbsforceerr_in), // input wire gt0_txprbsforceerr_in
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .gt0_txdata_in                  (gt0_txdata_in), // input wire [31:0] gt0_txdata_in
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .gt0_gthtxn_out                 (gt0_gthtxn_out), // output wire gt0_gthtxn_out
        .gt0_gthtxp_out                 (gt0_gthtxp_out), // output wire gt0_gthtxp_out
        //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        .gt0_txoutclk_out               (gt0_txoutclk_i), // output wire gt0_txoutclk_i
        .gt0_txoutclkfabric_out         (gt0_txoutclkfabric_out), // output wire gt0_txoutclkfabric_out
        .gt0_txoutclkpcs_out            (gt0_txoutclkpcs_out), // output wire gt0_txoutclkpcs_out
        //----------- Transmit Ports - TX Initialization and Reset Ports -----------
        .gt0_txresetdone_out            (gt0_txresetdone_i), // output wire gt0_txresetdone_i
        //---------------- Transmit Ports - pattern Generator Ports ----------------
        .gt0_txprbssel_in               (gt0_txprbssel_in), // input wire [2:0] gt0_txprbssel_in
        //--------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        .gt0_txcharisk_in               (gt0_txcharisk_in), // input wire [3:0] gt0_txcharisk_in


        .gt1_rxpmaresetdone_out         (gt1_rxpmaresetdone_i),
        .gt1_txpmaresetdone_out         (gt1_txpmaresetdone_i),
 
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GT1  (X1Y29)

        //-------------------------- Channel - DRP Ports  --------------------------
        .gt1_drpaddr_in                 (gt1_drpaddr_in), // input wire [8:0] gt1_drpaddr_in
        .gt1_drpclk_in                  (gt1_drpclk_in), // input wire gt1_drpclk_in
        .gt1_drpdi_in                   (gt1_drpdi_in), // input wire [15:0] gt1_drpdi_in
        .gt1_drpdo_out                  (gt1_drpdo_out), // output wire [15:0] gt1_drpdo_out
        .gt1_drpen_in                   (gt1_drpen_in), // input wire gt1_drpen_in
        .gt1_drprdy_out                 (gt1_drprdy_out), // output wire gt1_drprdy_out
        .gt1_drpwe_in                   (gt1_drpwe_in), // input wire gt1_drpwe_in
        //------------------- RX Initialization and Reset Ports --------------------
        .gt1_eyescanreset_in            (gt1_eyescanreset_in), // input wire gt1_eyescanreset_in
        .gt1_rxuserrdy_in               (gt1_rxuserrdy_i), // input wire gt1_rxuserrdy_i
        //------------------------ RX Margin Analysis Ports ------------------------
        .gt1_eyescandataerror_out       (gt1_eyescandataerror_out), // output wire gt1_eyescandataerror_out
        .gt1_eyescantrigger_in          (gt1_eyescantrigger_in), // input wire gt1_eyescantrigger_in
        //----------------- Receive Ports - Digital Monitor Ports ------------------
        .gt1_dmonitorout_out            (gt1_dmonitorout_out), // output wire [14:0] gt1_dmonitorout_out
        //---------------- Receive Ports - FPGA RX Interface Ports -----------------
        .gt1_rxusrclk_in                (gt1_rxusrclk_in), // input wire gt1_rxusrclk_in
        .gt1_rxusrclk2_in               (gt1_rxusrclk2_in), // input wire gt1_rxusrclk2_in
        //---------------- Receive Ports - FPGA RX interface Ports -----------------
        .gt1_rxdata_out                 (gt1_rxdata_out), // output wire [31:0] gt1_rxdata_out
        //----------------- Receive Ports - Pattern Checker Ports ------------------
        .gt1_rxprbserr_out              (gt1_rxprbserr_out), // output wire gt1_rxprbserr_out
        .gt1_rxprbssel_in               (gt1_rxprbssel_in), // input wire [2:0] gt1_rxprbssel_in
        //----------------- Receive Ports - Pattern Checker ports ------------------
        .gt1_rxprbscntreset_in          (gt1_rxprbscntreset_in), // input wire gt1_rxprbscntreset_in
        //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
        .gt1_rxdisperr_out              (gt1_rxdisperr_out), // output wire [3:0] gt1_rxdisperr_out
        .gt1_rxnotintable_out           (gt1_rxnotintable_out), // output wire [3:0] gt1_rxnotintable_out
        //---------------------- Receive Ports - RX AFE Ports ----------------------
        .gt1_gthrxn_in                  (gt1_gthrxn_in), // input wire gt1_gthrxn_in
        //------------ Receive Ports - RX Byte and Word Alignment Ports ------------
        .gt1_rxmcommaalignen_in         (gt1_rxmcommaalignen_in), // input wire gt1_rxmcommaalignen_in
        .gt1_rxpcommaalignen_in         (gt1_rxpcommaalignen_in), // input wire gt1_rxpcommaalignen_in
        //---------------- Receive Ports - RX Channel Bonding Ports ----------------
        .gt1_rxchanbondseq_out          (gt1_rxchanbondseq_out), // output wire gt1_rxchanbondseq_out
        .gt1_rxchbonden_in              (gt1_rxchbonden_in), // input wire gt1_rxchbonden_in
        .gt1_rxchbondlevel_in           (gt1_rxchbondlevel_in), // input wire [2:0] gt1_rxchbondlevel_in
        .gt1_rxchbondmaster_in          (gt1_rxchbondmaster_in), // input wire gt1_rxchbondmaster_in
        .gt1_rxchbondo_out              (gt1_rxchbondo_out), // output wire [4:0] gt1_rxchbondo_out
        .gt1_rxchbondslave_in           (gt1_rxchbondslave_in), // input wire gt1_rxchbondslave_in
        //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
        .gt1_rxchanisaligned_out        (gt1_rxchanisaligned_out), // output wire gt1_rxchanisaligned_out
        .gt1_rxchanrealign_out          (gt1_rxchanrealign_out), // output wire gt1_rxchanrealign_out
        //------------------- Receive Ports - RX Equalizer Ports -------------------
        .gt1_rxdfeagchold_in            (gt1_rxdfeagchold_i), // input wire gt1_rxdfeagchold_i
        .gt1_rxdfelfhold_in             (gt1_rxdfelfhold_i), // input wire gt1_rxdfelfhold_i
        .gt1_rxmonitorout_out           (gt1_rxmonitorout_out), // output wire [6:0] gt1_rxmonitorout_out
        .gt1_rxmonitorsel_in            (gt1_rxmonitorsel_in), // input wire [1:0] gt1_rxmonitorsel_in
        //------------- Receive Ports - RX Fabric Output Control Ports -------------
        .gt1_rxoutclk_out               (gt1_rxoutclk_i), // output wire gt1_rxoutclk_i
        //----------- Receive Ports - RX Initialization and Reset Ports ------------
        .gt1_gtrxreset_in               (gt1_gtrxreset_i), // input wire gt1_gtrxreset_i
        //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        .gt1_rxcharisk_out              (gt1_rxcharisk_out), // output wire [3:0] gt1_rxcharisk_out
        //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
        .gt1_rxchbondi_in               (gt1_rxchbondi_in), // input wire [4:0] gt1_rxchbondi_in
        //---------------------- Receive Ports -RX AFE Ports -----------------------
        .gt1_gthrxp_in                  (gt1_gthrxp_in), // input wire gt1_gthrxp_in
        //------------ Receive Ports -RX Initialization and Reset Ports ------------
        .gt1_rxresetdone_out            (gt1_rxresetdone_i), // output wire gt1_rxresetdone_i
        //------------------- TX Initialization and Reset Ports --------------------
        .gt1_gttxreset_in               (gt1_gttxreset_i), // input wire gt1_gttxreset_i
        .gt1_txuserrdy_in               (gt1_txuserrdy_i), // input wire gt1_txuserrdy_i
        //-------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        .gt1_txchardispmode_in          (gt1_txchardispmode_in), // input wire [3:0] gt1_txchardispmode_in
        .gt1_txchardispval_in           (gt1_txchardispval_in), // input wire [3:0] gt1_txchardispval_in
        //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
        .gt1_txusrclk_in                (gt1_txusrclk_in), // input wire gt1_txusrclk_in
        .gt1_txusrclk2_in               (gt1_txusrclk2_in), // input wire gt1_txusrclk2_in
        //---------------- Transmit Ports - Pattern Generator Ports ----------------
        .gt1_txprbsforceerr_in          (gt1_txprbsforceerr_in), // input wire gt1_txprbsforceerr_in
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .gt1_txdata_in                  (gt1_txdata_in), // input wire [31:0] gt1_txdata_in
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .gt1_gthtxn_out                 (gt1_gthtxn_out), // output wire gt1_gthtxn_out
        .gt1_gthtxp_out                 (gt1_gthtxp_out), // output wire gt1_gthtxp_out
        //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        .gt1_txoutclk_out               (gt1_txoutclk_i), // output wire gt1_txoutclk_i
        .gt1_txoutclkfabric_out         (gt1_txoutclkfabric_out), // output wire gt1_txoutclkfabric_out
        .gt1_txoutclkpcs_out            (gt1_txoutclkpcs_out), // output wire gt1_txoutclkpcs_out
        //----------- Transmit Ports - TX Initialization and Reset Ports -----------
        .gt1_txresetdone_out            (gt1_txresetdone_i), // output wire gt1_txresetdone_i
        //---------------- Transmit Ports - pattern Generator Ports ----------------
        .gt1_txprbssel_in               (gt1_txprbssel_in), // input wire [2:0] gt1_txprbssel_in
        //--------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        .gt1_txcharisk_in               (gt1_txcharisk_in), // input wire [3:0] gt1_txcharisk_in


        .gt2_rxpmaresetdone_out         (gt2_rxpmaresetdone_i),
        .gt2_txpmaresetdone_out         (gt2_txpmaresetdone_i),
 
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GT2  (X1Y32)

        //-------------------------- Channel - DRP Ports  --------------------------
        .gt2_drpaddr_in                 (gt2_drpaddr_in), // input wire [8:0] gt2_drpaddr_in
        .gt2_drpclk_in                  (gt2_drpclk_in), // input wire gt2_drpclk_in
        .gt2_drpdi_in                   (gt2_drpdi_in), // input wire [15:0] gt2_drpdi_in
        .gt2_drpdo_out                  (gt2_drpdo_out), // output wire [15:0] gt2_drpdo_out
        .gt2_drpen_in                   (gt2_drpen_in), // input wire gt2_drpen_in
        .gt2_drprdy_out                 (gt2_drprdy_out), // output wire gt2_drprdy_out
        .gt2_drpwe_in                   (gt2_drpwe_in), // input wire gt2_drpwe_in
        //------------------- RX Initialization and Reset Ports --------------------
        .gt2_eyescanreset_in            (gt2_eyescanreset_in), // input wire gt2_eyescanreset_in
        .gt2_rxuserrdy_in               (gt2_rxuserrdy_i), // input wire gt2_rxuserrdy_i
        //------------------------ RX Margin Analysis Ports ------------------------
        .gt2_eyescandataerror_out       (gt2_eyescandataerror_out), // output wire gt2_eyescandataerror_out
        .gt2_eyescantrigger_in          (gt2_eyescantrigger_in), // input wire gt2_eyescantrigger_in
        //----------------- Receive Ports - Digital Monitor Ports ------------------
        .gt2_dmonitorout_out            (gt2_dmonitorout_out), // output wire [14:0] gt2_dmonitorout_out
        //---------------- Receive Ports - FPGA RX Interface Ports -----------------
        .gt2_rxusrclk_in                (gt2_rxusrclk_in), // input wire gt2_rxusrclk_in
        .gt2_rxusrclk2_in               (gt2_rxusrclk2_in), // input wire gt2_rxusrclk2_in
        //---------------- Receive Ports - FPGA RX interface Ports -----------------
        .gt2_rxdata_out                 (gt2_rxdata_out), // output wire [31:0] gt2_rxdata_out
        //----------------- Receive Ports - Pattern Checker Ports ------------------
        .gt2_rxprbserr_out              (gt2_rxprbserr_out), // output wire gt2_rxprbserr_out
        .gt2_rxprbssel_in               (gt2_rxprbssel_in), // input wire [2:0] gt2_rxprbssel_in
        //----------------- Receive Ports - Pattern Checker ports ------------------
        .gt2_rxprbscntreset_in          (gt2_rxprbscntreset_in), // input wire gt2_rxprbscntreset_in
        //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
        .gt2_rxdisperr_out              (gt2_rxdisperr_out), // output wire [3:0] gt2_rxdisperr_out
        .gt2_rxnotintable_out           (gt2_rxnotintable_out), // output wire [3:0] gt2_rxnotintable_out
        //---------------------- Receive Ports - RX AFE Ports ----------------------
        .gt2_gthrxn_in                  (gt2_gthrxn_in), // input wire gt2_gthrxn_in
        //------------ Receive Ports - RX Byte and Word Alignment Ports ------------
        .gt2_rxmcommaalignen_in         (gt2_rxmcommaalignen_in), // input wire gt2_rxmcommaalignen_in
        .gt2_rxpcommaalignen_in         (gt2_rxpcommaalignen_in), // input wire gt2_rxpcommaalignen_in
        //---------------- Receive Ports - RX Channel Bonding Ports ----------------
        .gt2_rxchanbondseq_out          (gt2_rxchanbondseq_out), // output wire gt2_rxchanbondseq_out
        .gt2_rxchbonden_in              (gt2_rxchbonden_in), // input wire gt2_rxchbonden_in
        .gt2_rxchbondlevel_in           (gt2_rxchbondlevel_in), // input wire [2:0] gt2_rxchbondlevel_in
        .gt2_rxchbondmaster_in          (gt2_rxchbondmaster_in), // input wire gt2_rxchbondmaster_in
        .gt2_rxchbondo_out              (gt2_rxchbondo_out), // output wire [4:0] gt2_rxchbondo_out
        .gt2_rxchbondslave_in           (gt2_rxchbondslave_in), // input wire gt2_rxchbondslave_in
        //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
        .gt2_rxchanisaligned_out        (gt2_rxchanisaligned_out), // output wire gt2_rxchanisaligned_out
        .gt2_rxchanrealign_out          (gt2_rxchanrealign_out), // output wire gt2_rxchanrealign_out
        //------------------- Receive Ports - RX Equalizer Ports -------------------
        .gt2_rxdfeagchold_in            (gt2_rxdfeagchold_i), // input wire gt2_rxdfeagchold_i
        .gt2_rxdfelfhold_in             (gt2_rxdfelfhold_i), // input wire gt2_rxdfelfhold_i
        .gt2_rxmonitorout_out           (gt2_rxmonitorout_out), // output wire [6:0] gt2_rxmonitorout_out
        .gt2_rxmonitorsel_in            (gt2_rxmonitorsel_in), // input wire [1:0] gt2_rxmonitorsel_in
        //------------- Receive Ports - RX Fabric Output Control Ports -------------
        .gt2_rxoutclk_out               (gt2_rxoutclk_i), // output wire gt2_rxoutclk_i
        //----------- Receive Ports - RX Initialization and Reset Ports ------------
        .gt2_gtrxreset_in               (gt2_gtrxreset_i), // input wire gt2_gtrxreset_i
        //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        .gt2_rxcharisk_out              (gt2_rxcharisk_out), // output wire [3:0] gt2_rxcharisk_out
        //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
        .gt2_rxchbondi_in               (gt2_rxchbondi_in), // input wire [4:0] gt2_rxchbondi_in
        //---------------------- Receive Ports -RX AFE Ports -----------------------
        .gt2_gthrxp_in                  (gt2_gthrxp_in), // input wire gt2_gthrxp_in
        //------------ Receive Ports -RX Initialization and Reset Ports ------------
        .gt2_rxresetdone_out            (gt2_rxresetdone_i), // output wire gt2_rxresetdone_i
        //------------------- TX Initialization and Reset Ports --------------------
        .gt2_gttxreset_in               (gt2_gttxreset_i), // input wire gt2_gttxreset_i
        .gt2_txuserrdy_in               (gt2_txuserrdy_i), // input wire gt2_txuserrdy_i
        //-------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        .gt2_txchardispmode_in          (gt2_txchardispmode_in), // input wire [3:0] gt2_txchardispmode_in
        .gt2_txchardispval_in           (gt2_txchardispval_in), // input wire [3:0] gt2_txchardispval_in
        //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
        .gt2_txusrclk_in                (gt2_txusrclk_in), // input wire gt2_txusrclk_in
        .gt2_txusrclk2_in               (gt2_txusrclk2_in), // input wire gt2_txusrclk2_in
        //---------------- Transmit Ports - Pattern Generator Ports ----------------
        .gt2_txprbsforceerr_in          (gt2_txprbsforceerr_in), // input wire gt2_txprbsforceerr_in
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .gt2_txdata_in                  (gt2_txdata_in), // input wire [31:0] gt2_txdata_in
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .gt2_gthtxn_out                 (gt2_gthtxn_out), // output wire gt2_gthtxn_out
        .gt2_gthtxp_out                 (gt2_gthtxp_out), // output wire gt2_gthtxp_out
        //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        .gt2_txoutclk_out               (gt2_txoutclk_i), // output wire gt2_txoutclk_i
        .gt2_txoutclkfabric_out         (gt2_txoutclkfabric_out), // output wire gt2_txoutclkfabric_out
        .gt2_txoutclkpcs_out            (gt2_txoutclkpcs_out), // output wire gt2_txoutclkpcs_out
        //----------- Transmit Ports - TX Initialization and Reset Ports -----------
        .gt2_txresetdone_out            (gt2_txresetdone_i), // output wire gt2_txresetdone_i
        //---------------- Transmit Ports - pattern Generator Ports ----------------
        .gt2_txprbssel_in               (gt2_txprbssel_in), // input wire [2:0] gt2_txprbssel_in
        //--------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        .gt2_txcharisk_in               (gt2_txcharisk_in), // input wire [3:0] gt2_txcharisk_in


        .gt3_rxpmaresetdone_out         (gt3_rxpmaresetdone_i),
        .gt3_txpmaresetdone_out         (gt3_txpmaresetdone_i),
 
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GT3  (X1Y33)

        //-------------------------- Channel - DRP Ports  --------------------------
        .gt3_drpaddr_in                 (gt3_drpaddr_in), // input wire [8:0] gt3_drpaddr_in
        .gt3_drpclk_in                  (gt3_drpclk_in), // input wire gt3_drpclk_in
        .gt3_drpdi_in                   (gt3_drpdi_in), // input wire [15:0] gt3_drpdi_in
        .gt3_drpdo_out                  (gt3_drpdo_out), // output wire [15:0] gt3_drpdo_out
        .gt3_drpen_in                   (gt3_drpen_in), // input wire gt3_drpen_in
        .gt3_drprdy_out                 (gt3_drprdy_out), // output wire gt3_drprdy_out
        .gt3_drpwe_in                   (gt3_drpwe_in), // input wire gt3_drpwe_in
        //------------------- RX Initialization and Reset Ports --------------------
        .gt3_eyescanreset_in            (gt3_eyescanreset_in), // input wire gt3_eyescanreset_in
        .gt3_rxuserrdy_in               (gt3_rxuserrdy_i), // input wire gt3_rxuserrdy_i
        //------------------------ RX Margin Analysis Ports ------------------------
        .gt3_eyescandataerror_out       (gt3_eyescandataerror_out), // output wire gt3_eyescandataerror_out
        .gt3_eyescantrigger_in          (gt3_eyescantrigger_in), // input wire gt3_eyescantrigger_in
        //----------------- Receive Ports - Digital Monitor Ports ------------------
        .gt3_dmonitorout_out            (gt3_dmonitorout_out), // output wire [14:0] gt3_dmonitorout_out
        //---------------- Receive Ports - FPGA RX Interface Ports -----------------
        .gt3_rxusrclk_in                (gt3_rxusrclk_in), // input wire gt3_rxusrclk_in
        .gt3_rxusrclk2_in               (gt3_rxusrclk2_in), // input wire gt3_rxusrclk2_in
        //---------------- Receive Ports - FPGA RX interface Ports -----------------
        .gt3_rxdata_out                 (gt3_rxdata_out), // output wire [31:0] gt3_rxdata_out
        //----------------- Receive Ports - Pattern Checker Ports ------------------
        .gt3_rxprbserr_out              (gt3_rxprbserr_out), // output wire gt3_rxprbserr_out
        .gt3_rxprbssel_in               (gt3_rxprbssel_in), // input wire [2:0] gt3_rxprbssel_in
        //----------------- Receive Ports - Pattern Checker ports ------------------
        .gt3_rxprbscntreset_in          (gt3_rxprbscntreset_in), // input wire gt3_rxprbscntreset_in
        //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
        .gt3_rxdisperr_out              (gt3_rxdisperr_out), // output wire [3:0] gt3_rxdisperr_out
        .gt3_rxnotintable_out           (gt3_rxnotintable_out), // output wire [3:0] gt3_rxnotintable_out
        //---------------------- Receive Ports - RX AFE Ports ----------------------
        .gt3_gthrxn_in                  (gt3_gthrxn_in), // input wire gt3_gthrxn_in
        //------------ Receive Ports - RX Byte and Word Alignment Ports ------------
        .gt3_rxmcommaalignen_in         (gt3_rxmcommaalignen_in), // input wire gt3_rxmcommaalignen_in
        .gt3_rxpcommaalignen_in         (gt3_rxpcommaalignen_in), // input wire gt3_rxpcommaalignen_in
        //---------------- Receive Ports - RX Channel Bonding Ports ----------------
        .gt3_rxchanbondseq_out          (gt3_rxchanbondseq_out), // output wire gt3_rxchanbondseq_out
        .gt3_rxchbonden_in              (gt3_rxchbonden_in), // input wire gt3_rxchbonden_in
        .gt3_rxchbondlevel_in           (gt3_rxchbondlevel_in), // input wire [2:0] gt3_rxchbondlevel_in
        .gt3_rxchbondmaster_in          (gt3_rxchbondmaster_in), // input wire gt3_rxchbondmaster_in
        .gt3_rxchbondo_out              (gt3_rxchbondo_out), // output wire [4:0] gt3_rxchbondo_out
        .gt3_rxchbondslave_in           (gt3_rxchbondslave_in), // input wire gt3_rxchbondslave_in
        //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
        .gt3_rxchanisaligned_out        (gt3_rxchanisaligned_out), // output wire gt3_rxchanisaligned_out
        .gt3_rxchanrealign_out          (gt3_rxchanrealign_out), // output wire gt3_rxchanrealign_out
        //------------------- Receive Ports - RX Equalizer Ports -------------------
        .gt3_rxdfeagchold_in            (gt3_rxdfeagchold_i), // input wire gt3_rxdfeagchold_i
        .gt3_rxdfelfhold_in             (gt3_rxdfelfhold_i), // input wire gt3_rxdfelfhold_i
        .gt3_rxmonitorout_out           (gt3_rxmonitorout_out), // output wire [6:0] gt3_rxmonitorout_out
        .gt3_rxmonitorsel_in            (gt3_rxmonitorsel_in), // input wire [1:0] gt3_rxmonitorsel_in
        //------------- Receive Ports - RX Fabric Output Control Ports -------------
        .gt3_rxoutclk_out               (gt3_rxoutclk_i), // output wire gt3_rxoutclk_i
        //----------- Receive Ports - RX Initialization and Reset Ports ------------
        .gt3_gtrxreset_in               (gt3_gtrxreset_i), // input wire gt3_gtrxreset_i
        //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        .gt3_rxcharisk_out              (gt3_rxcharisk_out), // output wire [3:0] gt3_rxcharisk_out
        //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
        .gt3_rxchbondi_in               (gt3_rxchbondi_in), // input wire [4:0] gt3_rxchbondi_in
        //---------------------- Receive Ports -RX AFE Ports -----------------------
        .gt3_gthrxp_in                  (gt3_gthrxp_in), // input wire gt3_gthrxp_in
        //------------ Receive Ports -RX Initialization and Reset Ports ------------
        .gt3_rxresetdone_out            (gt3_rxresetdone_i), // output wire gt3_rxresetdone_i
        //------------------- TX Initialization and Reset Ports --------------------
        .gt3_gttxreset_in               (gt3_gttxreset_i), // input wire gt3_gttxreset_i
        .gt3_txuserrdy_in               (gt3_txuserrdy_i), // input wire gt3_txuserrdy_i
        //-------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        .gt3_txchardispmode_in          (gt3_txchardispmode_in), // input wire [3:0] gt3_txchardispmode_in
        .gt3_txchardispval_in           (gt3_txchardispval_in), // input wire [3:0] gt3_txchardispval_in
        //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
        .gt3_txusrclk_in                (gt3_txusrclk_in), // input wire gt3_txusrclk_in
        .gt3_txusrclk2_in               (gt3_txusrclk2_in), // input wire gt3_txusrclk2_in
        //---------------- Transmit Ports - Pattern Generator Ports ----------------
        .gt3_txprbsforceerr_in          (gt3_txprbsforceerr_in), // input wire gt3_txprbsforceerr_in
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .gt3_txdata_in                  (gt3_txdata_in), // input wire [31:0] gt3_txdata_in
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .gt3_gthtxn_out                 (gt3_gthtxn_out), // output wire gt3_gthtxn_out
        .gt3_gthtxp_out                 (gt3_gthtxp_out), // output wire gt3_gthtxp_out
        //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        .gt3_txoutclk_out               (gt3_txoutclk_i), // output wire gt3_txoutclk_i
        .gt3_txoutclkfabric_out         (gt3_txoutclkfabric_out), // output wire gt3_txoutclkfabric_out
        .gt3_txoutclkpcs_out            (gt3_txoutclkpcs_out), // output wire gt3_txoutclkpcs_out
        //----------- Transmit Ports - TX Initialization and Reset Ports -----------
        .gt3_txresetdone_out            (gt3_txresetdone_i), // output wire gt3_txresetdone_i
        //---------------- Transmit Ports - pattern Generator Ports ----------------
        .gt3_txprbssel_in               (gt3_txprbssel_in), // input wire [2:0] gt3_txprbssel_in
        //--------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        .gt3_txcharisk_in               (gt3_txcharisk_in), // input wire [3:0] gt3_txcharisk_in


        .gt4_rxpmaresetdone_out         (gt4_rxpmaresetdone_i),
        .gt4_txpmaresetdone_out         (gt4_txpmaresetdone_i),
 
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GT4  (X1Y34)

        //-------------------------- Channel - DRP Ports  --------------------------
        .gt4_drpaddr_in                 (gt4_drpaddr_in), // input wire [8:0] gt4_drpaddr_in
        .gt4_drpclk_in                  (gt4_drpclk_in), // input wire gt4_drpclk_in
        .gt4_drpdi_in                   (gt4_drpdi_in), // input wire [15:0] gt4_drpdi_in
        .gt4_drpdo_out                  (gt4_drpdo_out), // output wire [15:0] gt4_drpdo_out
        .gt4_drpen_in                   (gt4_drpen_in), // input wire gt4_drpen_in
        .gt4_drprdy_out                 (gt4_drprdy_out), // output wire gt4_drprdy_out
        .gt4_drpwe_in                   (gt4_drpwe_in), // input wire gt4_drpwe_in
        //------------------- RX Initialization and Reset Ports --------------------
        .gt4_eyescanreset_in            (gt4_eyescanreset_in), // input wire gt4_eyescanreset_in
        .gt4_rxuserrdy_in               (gt4_rxuserrdy_i), // input wire gt4_rxuserrdy_i
        //------------------------ RX Margin Analysis Ports ------------------------
        .gt4_eyescandataerror_out       (gt4_eyescandataerror_out), // output wire gt4_eyescandataerror_out
        .gt4_eyescantrigger_in          (gt4_eyescantrigger_in), // input wire gt4_eyescantrigger_in
        //----------------- Receive Ports - Digital Monitor Ports ------------------
        .gt4_dmonitorout_out            (gt4_dmonitorout_out), // output wire [14:0] gt4_dmonitorout_out
        //---------------- Receive Ports - FPGA RX Interface Ports -----------------
        .gt4_rxusrclk_in                (gt4_rxusrclk_in), // input wire gt4_rxusrclk_in
        .gt4_rxusrclk2_in               (gt4_rxusrclk2_in), // input wire gt4_rxusrclk2_in
        //---------------- Receive Ports - FPGA RX interface Ports -----------------
        .gt4_rxdata_out                 (gt4_rxdata_out), // output wire [31:0] gt4_rxdata_out
        //----------------- Receive Ports - Pattern Checker Ports ------------------
        .gt4_rxprbserr_out              (gt4_rxprbserr_out), // output wire gt4_rxprbserr_out
        .gt4_rxprbssel_in               (gt4_rxprbssel_in), // input wire [2:0] gt4_rxprbssel_in
        //----------------- Receive Ports - Pattern Checker ports ------------------
        .gt4_rxprbscntreset_in          (gt4_rxprbscntreset_in), // input wire gt4_rxprbscntreset_in
        //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
        .gt4_rxdisperr_out              (gt4_rxdisperr_out), // output wire [3:0] gt4_rxdisperr_out
        .gt4_rxnotintable_out           (gt4_rxnotintable_out), // output wire [3:0] gt4_rxnotintable_out
        //---------------------- Receive Ports - RX AFE Ports ----------------------
        .gt4_gthrxn_in                  (gt4_gthrxn_in), // input wire gt4_gthrxn_in
        //------------ Receive Ports - RX Byte and Word Alignment Ports ------------
        .gt4_rxmcommaalignen_in         (gt4_rxmcommaalignen_in), // input wire gt4_rxmcommaalignen_in
        .gt4_rxpcommaalignen_in         (gt4_rxpcommaalignen_in), // input wire gt4_rxpcommaalignen_in
        //---------------- Receive Ports - RX Channel Bonding Ports ----------------
        .gt4_rxchanbondseq_out          (gt4_rxchanbondseq_out), // output wire gt4_rxchanbondseq_out
        .gt4_rxchbonden_in              (gt4_rxchbonden_in), // input wire gt4_rxchbonden_in
        .gt4_rxchbondlevel_in           (gt4_rxchbondlevel_in), // input wire [2:0] gt4_rxchbondlevel_in
        .gt4_rxchbondmaster_in          (gt4_rxchbondmaster_in), // input wire gt4_rxchbondmaster_in
        .gt4_rxchbondo_out              (gt4_rxchbondo_out), // output wire [4:0] gt4_rxchbondo_out
        .gt4_rxchbondslave_in           (gt4_rxchbondslave_in), // input wire gt4_rxchbondslave_in
        //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
        .gt4_rxchanisaligned_out        (gt4_rxchanisaligned_out), // output wire gt4_rxchanisaligned_out
        .gt4_rxchanrealign_out          (gt4_rxchanrealign_out), // output wire gt4_rxchanrealign_out
        //------------------- Receive Ports - RX Equalizer Ports -------------------
        .gt4_rxdfeagchold_in            (gt4_rxdfeagchold_i), // input wire gt4_rxdfeagchold_i
        .gt4_rxdfelfhold_in             (gt4_rxdfelfhold_i), // input wire gt4_rxdfelfhold_i
        .gt4_rxmonitorout_out           (gt4_rxmonitorout_out), // output wire [6:0] gt4_rxmonitorout_out
        .gt4_rxmonitorsel_in            (gt4_rxmonitorsel_in), // input wire [1:0] gt4_rxmonitorsel_in
        //------------- Receive Ports - RX Fabric Output Control Ports -------------
        .gt4_rxoutclk_out               (gt4_rxoutclk_i), // output wire gt4_rxoutclk_i
        //----------- Receive Ports - RX Initialization and Reset Ports ------------
        .gt4_gtrxreset_in               (gt4_gtrxreset_i), // input wire gt4_gtrxreset_i
        //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        .gt4_rxcharisk_out              (gt4_rxcharisk_out), // output wire [3:0] gt4_rxcharisk_out
        //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
        .gt4_rxchbondi_in               (gt4_rxchbondi_in), // input wire [4:0] gt4_rxchbondi_in
        //---------------------- Receive Ports -RX AFE Ports -----------------------
        .gt4_gthrxp_in                  (gt4_gthrxp_in), // input wire gt4_gthrxp_in
        //------------ Receive Ports -RX Initialization and Reset Ports ------------
        .gt4_rxresetdone_out            (gt4_rxresetdone_i), // output wire gt4_rxresetdone_i
        //------------------- TX Initialization and Reset Ports --------------------
        .gt4_gttxreset_in               (gt4_gttxreset_i), // input wire gt4_gttxreset_i
        .gt4_txuserrdy_in               (gt4_txuserrdy_i), // input wire gt4_txuserrdy_i
        //-------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        .gt4_txchardispmode_in          (gt4_txchardispmode_in), // input wire [3:0] gt4_txchardispmode_in
        .gt4_txchardispval_in           (gt4_txchardispval_in), // input wire [3:0] gt4_txchardispval_in
        //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
        .gt4_txusrclk_in                (gt4_txusrclk_in), // input wire gt4_txusrclk_in
        .gt4_txusrclk2_in               (gt4_txusrclk2_in), // input wire gt4_txusrclk2_in
        //---------------- Transmit Ports - Pattern Generator Ports ----------------
        .gt4_txprbsforceerr_in          (gt4_txprbsforceerr_in), // input wire gt4_txprbsforceerr_in
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .gt4_txdata_in                  (gt4_txdata_in), // input wire [31:0] gt4_txdata_in
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .gt4_gthtxn_out                 (gt4_gthtxn_out), // output wire gt4_gthtxn_out
        .gt4_gthtxp_out                 (gt4_gthtxp_out), // output wire gt4_gthtxp_out
        //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        .gt4_txoutclk_out               (gt4_txoutclk_i), // output wire gt4_txoutclk_i
        .gt4_txoutclkfabric_out         (gt4_txoutclkfabric_out), // output wire gt4_txoutclkfabric_out
        .gt4_txoutclkpcs_out            (gt4_txoutclkpcs_out), // output wire gt4_txoutclkpcs_out
        //----------- Transmit Ports - TX Initialization and Reset Ports -----------
        .gt4_txresetdone_out            (gt4_txresetdone_i), // output wire gt4_txresetdone_i
        //---------------- Transmit Ports - pattern Generator Ports ----------------
        .gt4_txprbssel_in               (gt4_txprbssel_in), // input wire [2:0] gt4_txprbssel_in
        //--------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        .gt4_txcharisk_in               (gt4_txcharisk_in), // input wire [3:0] gt4_txcharisk_in


        .gt5_rxpmaresetdone_out         (gt5_rxpmaresetdone_i),
        .gt5_txpmaresetdone_out         (gt5_txpmaresetdone_i),
 
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GT5  (X1Y35)

        //-------------------------- Channel - DRP Ports  --------------------------
        .gt5_drpaddr_in                 (gt5_drpaddr_in), // input wire [8:0] gt5_drpaddr_in
        .gt5_drpclk_in                  (gt5_drpclk_in), // input wire gt5_drpclk_in
        .gt5_drpdi_in                   (gt5_drpdi_in), // input wire [15:0] gt5_drpdi_in
        .gt5_drpdo_out                  (gt5_drpdo_out), // output wire [15:0] gt5_drpdo_out
        .gt5_drpen_in                   (gt5_drpen_in), // input wire gt5_drpen_in
        .gt5_drprdy_out                 (gt5_drprdy_out), // output wire gt5_drprdy_out
        .gt5_drpwe_in                   (gt5_drpwe_in), // input wire gt5_drpwe_in
        //------------------- RX Initialization and Reset Ports --------------------
        .gt5_eyescanreset_in            (gt5_eyescanreset_in), // input wire gt5_eyescanreset_in
        .gt5_rxuserrdy_in               (gt5_rxuserrdy_i), // input wire gt5_rxuserrdy_i
        //------------------------ RX Margin Analysis Ports ------------------------
        .gt5_eyescandataerror_out       (gt5_eyescandataerror_out), // output wire gt5_eyescandataerror_out
        .gt5_eyescantrigger_in          (gt5_eyescantrigger_in), // input wire gt5_eyescantrigger_in
        //----------------- Receive Ports - Digital Monitor Ports ------------------
        .gt5_dmonitorout_out            (gt5_dmonitorout_out), // output wire [14:0] gt5_dmonitorout_out
        //---------------- Receive Ports - FPGA RX Interface Ports -----------------
        .gt5_rxusrclk_in                (gt5_rxusrclk_in), // input wire gt5_rxusrclk_in
        .gt5_rxusrclk2_in               (gt5_rxusrclk2_in), // input wire gt5_rxusrclk2_in
        //---------------- Receive Ports - FPGA RX interface Ports -----------------
        .gt5_rxdata_out                 (gt5_rxdata_out), // output wire [31:0] gt5_rxdata_out
        //----------------- Receive Ports - Pattern Checker Ports ------------------
        .gt5_rxprbserr_out              (gt5_rxprbserr_out), // output wire gt5_rxprbserr_out
        .gt5_rxprbssel_in               (gt5_rxprbssel_in), // input wire [2:0] gt5_rxprbssel_in
        //----------------- Receive Ports - Pattern Checker ports ------------------
        .gt5_rxprbscntreset_in          (gt5_rxprbscntreset_in), // input wire gt5_rxprbscntreset_in
        //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
        .gt5_rxdisperr_out              (gt5_rxdisperr_out), // output wire [3:0] gt5_rxdisperr_out
        .gt5_rxnotintable_out           (gt5_rxnotintable_out), // output wire [3:0] gt5_rxnotintable_out
        //---------------------- Receive Ports - RX AFE Ports ----------------------
        .gt5_gthrxn_in                  (gt5_gthrxn_in), // input wire gt5_gthrxn_in
        //------------ Receive Ports - RX Byte and Word Alignment Ports ------------
        .gt5_rxmcommaalignen_in         (gt5_rxmcommaalignen_in), // input wire gt5_rxmcommaalignen_in
        .gt5_rxpcommaalignen_in         (gt5_rxpcommaalignen_in), // input wire gt5_rxpcommaalignen_in
        //---------------- Receive Ports - RX Channel Bonding Ports ----------------
        .gt5_rxchanbondseq_out          (gt5_rxchanbondseq_out), // output wire gt5_rxchanbondseq_out
        .gt5_rxchbonden_in              (gt5_rxchbonden_in), // input wire gt5_rxchbonden_in
        .gt5_rxchbondlevel_in           (gt5_rxchbondlevel_in), // input wire [2:0] gt5_rxchbondlevel_in
        .gt5_rxchbondmaster_in          (gt5_rxchbondmaster_in), // input wire gt5_rxchbondmaster_in
        .gt5_rxchbondo_out              (gt5_rxchbondo_out), // output wire [4:0] gt5_rxchbondo_out
        .gt5_rxchbondslave_in           (gt5_rxchbondslave_in), // input wire gt5_rxchbondslave_in
        //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
        .gt5_rxchanisaligned_out        (gt5_rxchanisaligned_out), // output wire gt5_rxchanisaligned_out
        .gt5_rxchanrealign_out          (gt5_rxchanrealign_out), // output wire gt5_rxchanrealign_out
        //------------------- Receive Ports - RX Equalizer Ports -------------------
        .gt5_rxdfeagchold_in            (gt5_rxdfeagchold_i), // input wire gt5_rxdfeagchold_i
        .gt5_rxdfelfhold_in             (gt5_rxdfelfhold_i), // input wire gt5_rxdfelfhold_i
        .gt5_rxmonitorout_out           (gt5_rxmonitorout_out), // output wire [6:0] gt5_rxmonitorout_out
        .gt5_rxmonitorsel_in            (gt5_rxmonitorsel_in), // input wire [1:0] gt5_rxmonitorsel_in
        //------------- Receive Ports - RX Fabric Output Control Ports -------------
        .gt5_rxoutclk_out               (gt5_rxoutclk_i), // output wire gt5_rxoutclk_i
        //----------- Receive Ports - RX Initialization and Reset Ports ------------
        .gt5_gtrxreset_in               (gt5_gtrxreset_i), // input wire gt5_gtrxreset_i
        //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        .gt5_rxcharisk_out              (gt5_rxcharisk_out), // output wire [3:0] gt5_rxcharisk_out
        //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
        .gt5_rxchbondi_in               (gt5_rxchbondi_in), // input wire [4:0] gt5_rxchbondi_in
        //---------------------- Receive Ports -RX AFE Ports -----------------------
        .gt5_gthrxp_in                  (gt5_gthrxp_in), // input wire gt5_gthrxp_in
        //------------ Receive Ports -RX Initialization and Reset Ports ------------
        .gt5_rxresetdone_out            (gt5_rxresetdone_i), // output wire gt5_rxresetdone_i
        //------------------- TX Initialization and Reset Ports --------------------
        .gt5_gttxreset_in               (gt5_gttxreset_i), // input wire gt5_gttxreset_i
        .gt5_txuserrdy_in               (gt5_txuserrdy_i), // input wire gt5_txuserrdy_i
        //-------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        .gt5_txchardispmode_in          (gt5_txchardispmode_in), // input wire [3:0] gt5_txchardispmode_in
        .gt5_txchardispval_in           (gt5_txchardispval_in), // input wire [3:0] gt5_txchardispval_in
        //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
        .gt5_txusrclk_in                (gt5_txusrclk_in), // input wire gt5_txusrclk_in
        .gt5_txusrclk2_in               (gt5_txusrclk2_in), // input wire gt5_txusrclk2_in
        //---------------- Transmit Ports - Pattern Generator Ports ----------------
        .gt5_txprbsforceerr_in          (gt5_txprbsforceerr_in), // input wire gt5_txprbsforceerr_in
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .gt5_txdata_in                  (gt5_txdata_in), // input wire [31:0] gt5_txdata_in
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .gt5_gthtxn_out                 (gt5_gthtxn_out), // output wire gt5_gthtxn_out
        .gt5_gthtxp_out                 (gt5_gthtxp_out), // output wire gt5_gthtxp_out
        //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        .gt5_txoutclk_out               (gt5_txoutclk_i), // output wire gt5_txoutclk_i
        .gt5_txoutclkfabric_out         (gt5_txoutclkfabric_out), // output wire gt5_txoutclkfabric_out
        .gt5_txoutclkpcs_out            (gt5_txoutclkpcs_out), // output wire gt5_txoutclkpcs_out
        //----------- Transmit Ports - TX Initialization and Reset Ports -----------
        .gt5_txresetdone_out            (gt5_txresetdone_i), // output wire gt5_txresetdone_i
        //---------------- Transmit Ports - pattern Generator Ports ----------------
        .gt5_txprbssel_in               (gt5_txprbssel_in), // input wire [2:0] gt5_txprbssel_in
        //--------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        .gt5_txcharisk_in               (gt5_txcharisk_in), // input wire [3:0] gt5_txcharisk_in


        .gt6_rxpmaresetdone_out         (gt6_rxpmaresetdone_i),
        .gt6_txpmaresetdone_out         (gt6_txpmaresetdone_i),
 
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GT6  (X1Y36)

        //-------------------------- Channel - DRP Ports  --------------------------
        .gt6_drpaddr_in                 (gt6_drpaddr_in), // input wire [8:0] gt6_drpaddr_in
        .gt6_drpclk_in                  (gt6_drpclk_in), // input wire gt6_drpclk_in
        .gt6_drpdi_in                   (gt6_drpdi_in), // input wire [15:0] gt6_drpdi_in
        .gt6_drpdo_out                  (gt6_drpdo_out), // output wire [15:0] gt6_drpdo_out
        .gt6_drpen_in                   (gt6_drpen_in), // input wire gt6_drpen_in
        .gt6_drprdy_out                 (gt6_drprdy_out), // output wire gt6_drprdy_out
        .gt6_drpwe_in                   (gt6_drpwe_in), // input wire gt6_drpwe_in
        //------------------- RX Initialization and Reset Ports --------------------
        .gt6_eyescanreset_in            (gt6_eyescanreset_in), // input wire gt6_eyescanreset_in
        .gt6_rxuserrdy_in               (gt6_rxuserrdy_i), // input wire gt6_rxuserrdy_i
        //------------------------ RX Margin Analysis Ports ------------------------
        .gt6_eyescandataerror_out       (gt6_eyescandataerror_out), // output wire gt6_eyescandataerror_out
        .gt6_eyescantrigger_in          (gt6_eyescantrigger_in), // input wire gt6_eyescantrigger_in
        //----------------- Receive Ports - Digital Monitor Ports ------------------
        .gt6_dmonitorout_out            (gt6_dmonitorout_out), // output wire [14:0] gt6_dmonitorout_out
        //---------------- Receive Ports - FPGA RX Interface Ports -----------------
        .gt6_rxusrclk_in                (gt6_rxusrclk_in), // input wire gt6_rxusrclk_in
        .gt6_rxusrclk2_in               (gt6_rxusrclk2_in), // input wire gt6_rxusrclk2_in
        //---------------- Receive Ports - FPGA RX interface Ports -----------------
        .gt6_rxdata_out                 (gt6_rxdata_out), // output wire [31:0] gt6_rxdata_out
        //----------------- Receive Ports - Pattern Checker Ports ------------------
        .gt6_rxprbserr_out              (gt6_rxprbserr_out), // output wire gt6_rxprbserr_out
        .gt6_rxprbssel_in               (gt6_rxprbssel_in), // input wire [2:0] gt6_rxprbssel_in
        //----------------- Receive Ports - Pattern Checker ports ------------------
        .gt6_rxprbscntreset_in          (gt6_rxprbscntreset_in), // input wire gt6_rxprbscntreset_in
        //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
        .gt6_rxdisperr_out              (gt6_rxdisperr_out), // output wire [3:0] gt6_rxdisperr_out
        .gt6_rxnotintable_out           (gt6_rxnotintable_out), // output wire [3:0] gt6_rxnotintable_out
        //---------------------- Receive Ports - RX AFE Ports ----------------------
        .gt6_gthrxn_in                  (gt6_gthrxn_in), // input wire gt6_gthrxn_in
        //------------ Receive Ports - RX Byte and Word Alignment Ports ------------
        .gt6_rxmcommaalignen_in         (gt6_rxmcommaalignen_in), // input wire gt6_rxmcommaalignen_in
        .gt6_rxpcommaalignen_in         (gt6_rxpcommaalignen_in), // input wire gt6_rxpcommaalignen_in
        //---------------- Receive Ports - RX Channel Bonding Ports ----------------
        .gt6_rxchanbondseq_out          (gt6_rxchanbondseq_out), // output wire gt6_rxchanbondseq_out
        .gt6_rxchbonden_in              (gt6_rxchbonden_in), // input wire gt6_rxchbonden_in
        .gt6_rxchbondlevel_in           (gt6_rxchbondlevel_in), // input wire [2:0] gt6_rxchbondlevel_in
        .gt6_rxchbondmaster_in          (gt6_rxchbondmaster_in), // input wire gt6_rxchbondmaster_in
        .gt6_rxchbondo_out              (gt6_rxchbondo_out), // output wire [4:0] gt6_rxchbondo_out
        .gt6_rxchbondslave_in           (gt6_rxchbondslave_in), // input wire gt6_rxchbondslave_in
        //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
        .gt6_rxchanisaligned_out        (gt6_rxchanisaligned_out), // output wire gt6_rxchanisaligned_out
        .gt6_rxchanrealign_out          (gt6_rxchanrealign_out), // output wire gt6_rxchanrealign_out
        //------------------- Receive Ports - RX Equalizer Ports -------------------
        .gt6_rxdfeagchold_in            (gt6_rxdfeagchold_i), // input wire gt6_rxdfeagchold_i
        .gt6_rxdfelfhold_in             (gt6_rxdfelfhold_i), // input wire gt6_rxdfelfhold_i
        .gt6_rxmonitorout_out           (gt6_rxmonitorout_out), // output wire [6:0] gt6_rxmonitorout_out
        .gt6_rxmonitorsel_in            (gt6_rxmonitorsel_in), // input wire [1:0] gt6_rxmonitorsel_in
        //------------- Receive Ports - RX Fabric Output Control Ports -------------
        .gt6_rxoutclk_out               (gt6_rxoutclk_i), // output wire gt6_rxoutclk_i
        //----------- Receive Ports - RX Initialization and Reset Ports ------------
        .gt6_gtrxreset_in               (gt6_gtrxreset_i), // input wire gt6_gtrxreset_i
        //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        .gt6_rxcharisk_out              (gt6_rxcharisk_out), // output wire [3:0] gt6_rxcharisk_out
        //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
        .gt6_rxchbondi_in               (gt6_rxchbondi_in), // input wire [4:0] gt6_rxchbondi_in
        //---------------------- Receive Ports -RX AFE Ports -----------------------
        .gt6_gthrxp_in                  (gt6_gthrxp_in), // input wire gt6_gthrxp_in
        //------------ Receive Ports -RX Initialization and Reset Ports ------------
        .gt6_rxresetdone_out            (gt6_rxresetdone_i), // output wire gt6_rxresetdone_i
        //------------------- TX Initialization and Reset Ports --------------------
        .gt6_gttxreset_in               (gt6_gttxreset_i), // input wire gt6_gttxreset_i
        .gt6_txuserrdy_in               (gt6_txuserrdy_i), // input wire gt6_txuserrdy_i
        //-------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        .gt6_txchardispmode_in          (gt6_txchardispmode_in), // input wire [3:0] gt6_txchardispmode_in
        .gt6_txchardispval_in           (gt6_txchardispval_in), // input wire [3:0] gt6_txchardispval_in
        //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
        .gt6_txusrclk_in                (gt6_txusrclk_in), // input wire gt6_txusrclk_in
        .gt6_txusrclk2_in               (gt6_txusrclk2_in), // input wire gt6_txusrclk2_in
        //---------------- Transmit Ports - Pattern Generator Ports ----------------
        .gt6_txprbsforceerr_in          (gt6_txprbsforceerr_in), // input wire gt6_txprbsforceerr_in
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .gt6_txdata_in                  (gt6_txdata_in), // input wire [31:0] gt6_txdata_in
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .gt6_gthtxn_out                 (gt6_gthtxn_out), // output wire gt6_gthtxn_out
        .gt6_gthtxp_out                 (gt6_gthtxp_out), // output wire gt6_gthtxp_out
        //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        .gt6_txoutclk_out               (gt6_txoutclk_i), // output wire gt6_txoutclk_i
        .gt6_txoutclkfabric_out         (gt6_txoutclkfabric_out), // output wire gt6_txoutclkfabric_out
        .gt6_txoutclkpcs_out            (gt6_txoutclkpcs_out), // output wire gt6_txoutclkpcs_out
        //----------- Transmit Ports - TX Initialization and Reset Ports -----------
        .gt6_txresetdone_out            (gt6_txresetdone_i), // output wire gt6_txresetdone_i
        //---------------- Transmit Ports - pattern Generator Ports ----------------
        .gt6_txprbssel_in               (gt6_txprbssel_in), // input wire [2:0] gt6_txprbssel_in
        //--------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        .gt6_txcharisk_in               (gt6_txcharisk_in), // input wire [3:0] gt6_txcharisk_in


        .gt7_rxpmaresetdone_out         (gt7_rxpmaresetdone_i),
        .gt7_txpmaresetdone_out         (gt7_txpmaresetdone_i),
 
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GT7  (X1Y37)

        //-------------------------- Channel - DRP Ports  --------------------------
        .gt7_drpaddr_in                 (gt7_drpaddr_in), // input wire [8:0] gt7_drpaddr_in
        .gt7_drpclk_in                  (gt7_drpclk_in), // input wire gt7_drpclk_in
        .gt7_drpdi_in                   (gt7_drpdi_in), // input wire [15:0] gt7_drpdi_in
        .gt7_drpdo_out                  (gt7_drpdo_out), // output wire [15:0] gt7_drpdo_out
        .gt7_drpen_in                   (gt7_drpen_in), // input wire gt7_drpen_in
        .gt7_drprdy_out                 (gt7_drprdy_out), // output wire gt7_drprdy_out
        .gt7_drpwe_in                   (gt7_drpwe_in), // input wire gt7_drpwe_in
        //------------------- RX Initialization and Reset Ports --------------------
        .gt7_eyescanreset_in            (gt7_eyescanreset_in), // input wire gt7_eyescanreset_in
        .gt7_rxuserrdy_in               (gt7_rxuserrdy_i), // input wire gt7_rxuserrdy_i
        //------------------------ RX Margin Analysis Ports ------------------------
        .gt7_eyescandataerror_out       (gt7_eyescandataerror_out), // output wire gt7_eyescandataerror_out
        .gt7_eyescantrigger_in          (gt7_eyescantrigger_in), // input wire gt7_eyescantrigger_in
        //----------------- Receive Ports - Digital Monitor Ports ------------------
        .gt7_dmonitorout_out            (gt7_dmonitorout_out), // output wire [14:0] gt7_dmonitorout_out
        //---------------- Receive Ports - FPGA RX Interface Ports -----------------
        .gt7_rxusrclk_in                (gt7_rxusrclk_in), // input wire gt7_rxusrclk_in
        .gt7_rxusrclk2_in               (gt7_rxusrclk2_in), // input wire gt7_rxusrclk2_in
        //---------------- Receive Ports - FPGA RX interface Ports -----------------
        .gt7_rxdata_out                 (gt7_rxdata_out), // output wire [31:0] gt7_rxdata_out
        //----------------- Receive Ports - Pattern Checker Ports ------------------
        .gt7_rxprbserr_out              (gt7_rxprbserr_out), // output wire gt7_rxprbserr_out
        .gt7_rxprbssel_in               (gt7_rxprbssel_in), // input wire [2:0] gt7_rxprbssel_in
        //----------------- Receive Ports - Pattern Checker ports ------------------
        .gt7_rxprbscntreset_in          (gt7_rxprbscntreset_in), // input wire gt7_rxprbscntreset_in
        //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
        .gt7_rxdisperr_out              (gt7_rxdisperr_out), // output wire [3:0] gt7_rxdisperr_out
        .gt7_rxnotintable_out           (gt7_rxnotintable_out), // output wire [3:0] gt7_rxnotintable_out
        //---------------------- Receive Ports - RX AFE Ports ----------------------
        .gt7_gthrxn_in                  (gt7_gthrxn_in), // input wire gt7_gthrxn_in
        //------------ Receive Ports - RX Byte and Word Alignment Ports ------------
        .gt7_rxmcommaalignen_in         (gt7_rxmcommaalignen_in), // input wire gt7_rxmcommaalignen_in
        .gt7_rxpcommaalignen_in         (gt7_rxpcommaalignen_in), // input wire gt7_rxpcommaalignen_in
        //---------------- Receive Ports - RX Channel Bonding Ports ----------------
        .gt7_rxchanbondseq_out          (gt7_rxchanbondseq_out), // output wire gt7_rxchanbondseq_out
        .gt7_rxchbonden_in              (gt7_rxchbonden_in), // input wire gt7_rxchbonden_in
        .gt7_rxchbondlevel_in           (gt7_rxchbondlevel_in), // input wire [2:0] gt7_rxchbondlevel_in
        .gt7_rxchbondmaster_in          (gt7_rxchbondmaster_in), // input wire gt7_rxchbondmaster_in
        .gt7_rxchbondo_out              (gt7_rxchbondo_out), // output wire [4:0] gt7_rxchbondo_out
        .gt7_rxchbondslave_in           (gt7_rxchbondslave_in), // input wire gt7_rxchbondslave_in
        //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
        .gt7_rxchanisaligned_out        (gt7_rxchanisaligned_out), // output wire gt7_rxchanisaligned_out
        .gt7_rxchanrealign_out          (gt7_rxchanrealign_out), // output wire gt7_rxchanrealign_out
        //------------------- Receive Ports - RX Equalizer Ports -------------------
        .gt7_rxdfeagchold_in            (gt7_rxdfeagchold_i), // input wire gt7_rxdfeagchold_i
        .gt7_rxdfelfhold_in             (gt7_rxdfelfhold_i), // input wire gt7_rxdfelfhold_i
        .gt7_rxmonitorout_out           (gt7_rxmonitorout_out), // output wire [6:0] gt7_rxmonitorout_out
        .gt7_rxmonitorsel_in            (gt7_rxmonitorsel_in), // input wire [1:0] gt7_rxmonitorsel_in
        //------------- Receive Ports - RX Fabric Output Control Ports -------------
        .gt7_rxoutclk_out               (gt7_rxoutclk_i), // output wire gt7_rxoutclk_i
        //----------- Receive Ports - RX Initialization and Reset Ports ------------
        .gt7_gtrxreset_in               (gt7_gtrxreset_i), // input wire gt7_gtrxreset_i
        //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        .gt7_rxcharisk_out              (gt7_rxcharisk_out), // output wire [3:0] gt7_rxcharisk_out
        //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
        .gt7_rxchbondi_in               (gt7_rxchbondi_in), // input wire [4:0] gt7_rxchbondi_in
        //---------------------- Receive Ports -RX AFE Ports -----------------------
        .gt7_gthrxp_in                  (gt7_gthrxp_in), // input wire gt7_gthrxp_in
        //------------ Receive Ports -RX Initialization and Reset Ports ------------
        .gt7_rxresetdone_out            (gt7_rxresetdone_i), // output wire gt7_rxresetdone_i
        //------------------- TX Initialization and Reset Ports --------------------
        .gt7_gttxreset_in               (gt7_gttxreset_i), // input wire gt7_gttxreset_i
        .gt7_txuserrdy_in               (gt7_txuserrdy_i), // input wire gt7_txuserrdy_i
        //-------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        .gt7_txchardispmode_in          (gt7_txchardispmode_in), // input wire [3:0] gt7_txchardispmode_in
        .gt7_txchardispval_in           (gt7_txchardispval_in), // input wire [3:0] gt7_txchardispval_in
        //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
        .gt7_txusrclk_in                (gt7_txusrclk_in), // input wire gt7_txusrclk_in
        .gt7_txusrclk2_in               (gt7_txusrclk2_in), // input wire gt7_txusrclk2_in
        //---------------- Transmit Ports - Pattern Generator Ports ----------------
        .gt7_txprbsforceerr_in          (gt7_txprbsforceerr_in), // input wire gt7_txprbsforceerr_in
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .gt7_txdata_in                  (gt7_txdata_in), // input wire [31:0] gt7_txdata_in
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .gt7_gthtxn_out                 (gt7_gthtxn_out), // output wire gt7_gthtxn_out
        .gt7_gthtxp_out                 (gt7_gthtxp_out), // output wire gt7_gthtxp_out
        //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        .gt7_txoutclk_out               (gt7_txoutclk_i), // output wire gt7_txoutclk_i
        .gt7_txoutclkfabric_out         (gt7_txoutclkfabric_out), // output wire gt7_txoutclkfabric_out
        .gt7_txoutclkpcs_out            (gt7_txoutclkpcs_out), // output wire gt7_txoutclkpcs_out
        //----------- Transmit Ports - TX Initialization and Reset Ports -----------
        .gt7_txresetdone_out            (gt7_txresetdone_i), // output wire gt7_txresetdone_i
        //---------------- Transmit Ports - pattern Generator Ports ----------------
        .gt7_txprbssel_in               (gt7_txprbssel_in), // input wire [2:0] gt7_txprbssel_in
        //--------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        .gt7_txcharisk_in               (gt7_txcharisk_in), // input wire [3:0] gt7_txcharisk_in


        .gt8_rxpmaresetdone_out         (gt8_rxpmaresetdone_i),
        .gt8_txpmaresetdone_out         (gt8_txpmaresetdone_i),
 
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GT8  (X1Y38)

        //-------------------------- Channel - DRP Ports  --------------------------
        .gt8_drpaddr_in                 (gt8_drpaddr_in), // input wire [8:0] gt8_drpaddr_in
        .gt8_drpclk_in                  (gt8_drpclk_in), // input wire gt8_drpclk_in
        .gt8_drpdi_in                   (gt8_drpdi_in), // input wire [15:0] gt8_drpdi_in
        .gt8_drpdo_out                  (gt8_drpdo_out), // output wire [15:0] gt8_drpdo_out
        .gt8_drpen_in                   (gt8_drpen_in), // input wire gt8_drpen_in
        .gt8_drprdy_out                 (gt8_drprdy_out), // output wire gt8_drprdy_out
        .gt8_drpwe_in                   (gt8_drpwe_in), // input wire gt8_drpwe_in
        //------------------- RX Initialization and Reset Ports --------------------
        .gt8_eyescanreset_in            (gt8_eyescanreset_in), // input wire gt8_eyescanreset_in
        .gt8_rxuserrdy_in               (gt8_rxuserrdy_i), // input wire gt8_rxuserrdy_i
        //------------------------ RX Margin Analysis Ports ------------------------
        .gt8_eyescandataerror_out       (gt8_eyescandataerror_out), // output wire gt8_eyescandataerror_out
        .gt8_eyescantrigger_in          (gt8_eyescantrigger_in), // input wire gt8_eyescantrigger_in
        //----------------- Receive Ports - Digital Monitor Ports ------------------
        .gt8_dmonitorout_out            (gt8_dmonitorout_out), // output wire [14:0] gt8_dmonitorout_out
        //---------------- Receive Ports - FPGA RX Interface Ports -----------------
        .gt8_rxusrclk_in                (gt8_rxusrclk_in), // input wire gt8_rxusrclk_in
        .gt8_rxusrclk2_in               (gt8_rxusrclk2_in), // input wire gt8_rxusrclk2_in
        //---------------- Receive Ports - FPGA RX interface Ports -----------------
        .gt8_rxdata_out                 (gt8_rxdata_out), // output wire [31:0] gt8_rxdata_out
        //----------------- Receive Ports - Pattern Checker Ports ------------------
        .gt8_rxprbserr_out              (gt8_rxprbserr_out), // output wire gt8_rxprbserr_out
        .gt8_rxprbssel_in               (gt8_rxprbssel_in), // input wire [2:0] gt8_rxprbssel_in
        //----------------- Receive Ports - Pattern Checker ports ------------------
        .gt8_rxprbscntreset_in          (gt8_rxprbscntreset_in), // input wire gt8_rxprbscntreset_in
        //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
        .gt8_rxdisperr_out              (gt8_rxdisperr_out), // output wire [3:0] gt8_rxdisperr_out
        .gt8_rxnotintable_out           (gt8_rxnotintable_out), // output wire [3:0] gt8_rxnotintable_out
        //---------------------- Receive Ports - RX AFE Ports ----------------------
        .gt8_gthrxn_in                  (gt8_gthrxn_in), // input wire gt8_gthrxn_in
        //------------ Receive Ports - RX Byte and Word Alignment Ports ------------
        .gt8_rxmcommaalignen_in         (gt8_rxmcommaalignen_in), // input wire gt8_rxmcommaalignen_in
        .gt8_rxpcommaalignen_in         (gt8_rxpcommaalignen_in), // input wire gt8_rxpcommaalignen_in
        //---------------- Receive Ports - RX Channel Bonding Ports ----------------
        .gt8_rxchanbondseq_out          (gt8_rxchanbondseq_out), // output wire gt8_rxchanbondseq_out
        .gt8_rxchbonden_in              (gt8_rxchbonden_in), // input wire gt8_rxchbonden_in
        .gt8_rxchbondlevel_in           (gt8_rxchbondlevel_in), // input wire [2:0] gt8_rxchbondlevel_in
        .gt8_rxchbondmaster_in          (gt8_rxchbondmaster_in), // input wire gt8_rxchbondmaster_in
        .gt8_rxchbondo_out              (gt8_rxchbondo_out), // output wire [4:0] gt8_rxchbondo_out
        .gt8_rxchbondslave_in           (gt8_rxchbondslave_in), // input wire gt8_rxchbondslave_in
        //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
        .gt8_rxchanisaligned_out        (gt8_rxchanisaligned_out), // output wire gt8_rxchanisaligned_out
        .gt8_rxchanrealign_out          (gt8_rxchanrealign_out), // output wire gt8_rxchanrealign_out
        //------------------- Receive Ports - RX Equalizer Ports -------------------
        .gt8_rxdfeagchold_in            (gt8_rxdfeagchold_i), // input wire gt8_rxdfeagchold_i
        .gt8_rxdfelfhold_in             (gt8_rxdfelfhold_i), // input wire gt8_rxdfelfhold_i
        .gt8_rxmonitorout_out           (gt8_rxmonitorout_out), // output wire [6:0] gt8_rxmonitorout_out
        .gt8_rxmonitorsel_in            (gt8_rxmonitorsel_in), // input wire [1:0] gt8_rxmonitorsel_in
        //------------- Receive Ports - RX Fabric Output Control Ports -------------
        .gt8_rxoutclk_out               (gt8_rxoutclk_i), // output wire gt8_rxoutclk_i
        //----------- Receive Ports - RX Initialization and Reset Ports ------------
        .gt8_gtrxreset_in               (gt8_gtrxreset_i), // input wire gt8_gtrxreset_i
        //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        .gt8_rxcharisk_out              (gt8_rxcharisk_out), // output wire [3:0] gt8_rxcharisk_out
        //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
        .gt8_rxchbondi_in               (gt8_rxchbondi_in), // input wire [4:0] gt8_rxchbondi_in
        //---------------------- Receive Ports -RX AFE Ports -----------------------
        .gt8_gthrxp_in                  (gt8_gthrxp_in), // input wire gt8_gthrxp_in
        //------------ Receive Ports -RX Initialization and Reset Ports ------------
        .gt8_rxresetdone_out            (gt8_rxresetdone_i), // output wire gt8_rxresetdone_i
        //------------------- TX Initialization and Reset Ports --------------------
        .gt8_gttxreset_in               (gt8_gttxreset_i), // input wire gt8_gttxreset_i
        .gt8_txuserrdy_in               (gt8_txuserrdy_i), // input wire gt8_txuserrdy_i
        //-------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        .gt8_txchardispmode_in          (gt8_txchardispmode_in), // input wire [3:0] gt8_txchardispmode_in
        .gt8_txchardispval_in           (gt8_txchardispval_in), // input wire [3:0] gt8_txchardispval_in
        //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
        .gt8_txusrclk_in                (gt8_txusrclk_in), // input wire gt8_txusrclk_in
        .gt8_txusrclk2_in               (gt8_txusrclk2_in), // input wire gt8_txusrclk2_in
        //---------------- Transmit Ports - Pattern Generator Ports ----------------
        .gt8_txprbsforceerr_in          (gt8_txprbsforceerr_in), // input wire gt8_txprbsforceerr_in
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .gt8_txdata_in                  (gt8_txdata_in), // input wire [31:0] gt8_txdata_in
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .gt8_gthtxn_out                 (gt8_gthtxn_out), // output wire gt8_gthtxn_out
        .gt8_gthtxp_out                 (gt8_gthtxp_out), // output wire gt8_gthtxp_out
        //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        .gt8_txoutclk_out               (gt8_txoutclk_i), // output wire gt8_txoutclk_i
        .gt8_txoutclkfabric_out         (gt8_txoutclkfabric_out), // output wire gt8_txoutclkfabric_out
        .gt8_txoutclkpcs_out            (gt8_txoutclkpcs_out), // output wire gt8_txoutclkpcs_out
        //----------- Transmit Ports - TX Initialization and Reset Ports -----------
        .gt8_txresetdone_out            (gt8_txresetdone_i), // output wire gt8_txresetdone_i
        //---------------- Transmit Ports - pattern Generator Ports ----------------
        .gt8_txprbssel_in               (gt8_txprbssel_in), // input wire [2:0] gt8_txprbssel_in
        //--------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        .gt8_txcharisk_in               (gt8_txcharisk_in), // input wire [3:0] gt8_txcharisk_in


        .gt9_rxpmaresetdone_out         (gt9_rxpmaresetdone_i),
        .gt9_txpmaresetdone_out         (gt9_txpmaresetdone_i),
 
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GT9  (X1Y39)

        //-------------------------- Channel - DRP Ports  --------------------------
        .gt9_drpaddr_in                 (gt9_drpaddr_in), // input wire [8:0] gt9_drpaddr_in
        .gt9_drpclk_in                  (gt9_drpclk_in), // input wire gt9_drpclk_in
        .gt9_drpdi_in                   (gt9_drpdi_in), // input wire [15:0] gt9_drpdi_in
        .gt9_drpdo_out                  (gt9_drpdo_out), // output wire [15:0] gt9_drpdo_out
        .gt9_drpen_in                   (gt9_drpen_in), // input wire gt9_drpen_in
        .gt9_drprdy_out                 (gt9_drprdy_out), // output wire gt9_drprdy_out
        .gt9_drpwe_in                   (gt9_drpwe_in), // input wire gt9_drpwe_in
        //------------------- RX Initialization and Reset Ports --------------------
        .gt9_eyescanreset_in            (gt9_eyescanreset_in), // input wire gt9_eyescanreset_in
        .gt9_rxuserrdy_in               (gt9_rxuserrdy_i), // input wire gt9_rxuserrdy_i
        //------------------------ RX Margin Analysis Ports ------------------------
        .gt9_eyescandataerror_out       (gt9_eyescandataerror_out), // output wire gt9_eyescandataerror_out
        .gt9_eyescantrigger_in          (gt9_eyescantrigger_in), // input wire gt9_eyescantrigger_in
        //----------------- Receive Ports - Digital Monitor Ports ------------------
        .gt9_dmonitorout_out            (gt9_dmonitorout_out), // output wire [14:0] gt9_dmonitorout_out
        //---------------- Receive Ports - FPGA RX Interface Ports -----------------
        .gt9_rxusrclk_in                (gt9_rxusrclk_in), // input wire gt9_rxusrclk_in
        .gt9_rxusrclk2_in               (gt9_rxusrclk2_in), // input wire gt9_rxusrclk2_in
        //---------------- Receive Ports - FPGA RX interface Ports -----------------
        .gt9_rxdata_out                 (gt9_rxdata_out), // output wire [31:0] gt9_rxdata_out
        //----------------- Receive Ports - Pattern Checker Ports ------------------
        .gt9_rxprbserr_out              (gt9_rxprbserr_out), // output wire gt9_rxprbserr_out
        .gt9_rxprbssel_in               (gt9_rxprbssel_in), // input wire [2:0] gt9_rxprbssel_in
        //----------------- Receive Ports - Pattern Checker ports ------------------
        .gt9_rxprbscntreset_in          (gt9_rxprbscntreset_in), // input wire gt9_rxprbscntreset_in
        //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
        .gt9_rxdisperr_out              (gt9_rxdisperr_out), // output wire [3:0] gt9_rxdisperr_out
        .gt9_rxnotintable_out           (gt9_rxnotintable_out), // output wire [3:0] gt9_rxnotintable_out
        //---------------------- Receive Ports - RX AFE Ports ----------------------
        .gt9_gthrxn_in                  (gt9_gthrxn_in), // input wire gt9_gthrxn_in
        //------------ Receive Ports - RX Byte and Word Alignment Ports ------------
        .gt9_rxmcommaalignen_in         (gt9_rxmcommaalignen_in), // input wire gt9_rxmcommaalignen_in
        .gt9_rxpcommaalignen_in         (gt9_rxpcommaalignen_in), // input wire gt9_rxpcommaalignen_in
        //---------------- Receive Ports - RX Channel Bonding Ports ----------------
        .gt9_rxchanbondseq_out          (gt9_rxchanbondseq_out), // output wire gt9_rxchanbondseq_out
        .gt9_rxchbonden_in              (gt9_rxchbonden_in), // input wire gt9_rxchbonden_in
        .gt9_rxchbondlevel_in           (gt9_rxchbondlevel_in), // input wire [2:0] gt9_rxchbondlevel_in
        .gt9_rxchbondmaster_in          (gt9_rxchbondmaster_in), // input wire gt9_rxchbondmaster_in
        .gt9_rxchbondo_out              (gt9_rxchbondo_out), // output wire [4:0] gt9_rxchbondo_out
        .gt9_rxchbondslave_in           (gt9_rxchbondslave_in), // input wire gt9_rxchbondslave_in
        //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
        .gt9_rxchanisaligned_out        (gt9_rxchanisaligned_out), // output wire gt9_rxchanisaligned_out
        .gt9_rxchanrealign_out          (gt9_rxchanrealign_out), // output wire gt9_rxchanrealign_out
        //------------------- Receive Ports - RX Equalizer Ports -------------------
        .gt9_rxdfeagchold_in            (gt9_rxdfeagchold_i), // input wire gt9_rxdfeagchold_i
        .gt9_rxdfelfhold_in             (gt9_rxdfelfhold_i), // input wire gt9_rxdfelfhold_i
        .gt9_rxmonitorout_out           (gt9_rxmonitorout_out), // output wire [6:0] gt9_rxmonitorout_out
        .gt9_rxmonitorsel_in            (gt9_rxmonitorsel_in), // input wire [1:0] gt9_rxmonitorsel_in
        //------------- Receive Ports - RX Fabric Output Control Ports -------------
        .gt9_rxoutclk_out               (gt9_rxoutclk_i), // output wire gt9_rxoutclk_i
        //----------- Receive Ports - RX Initialization and Reset Ports ------------
        .gt9_gtrxreset_in               (gt9_gtrxreset_i), // input wire gt9_gtrxreset_i
        //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        .gt9_rxcharisk_out              (gt9_rxcharisk_out), // output wire [3:0] gt9_rxcharisk_out
        //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
        .gt9_rxchbondi_in               (gt9_rxchbondi_in), // input wire [4:0] gt9_rxchbondi_in
        //---------------------- Receive Ports -RX AFE Ports -----------------------
        .gt9_gthrxp_in                  (gt9_gthrxp_in), // input wire gt9_gthrxp_in
        //------------ Receive Ports -RX Initialization and Reset Ports ------------
        .gt9_rxresetdone_out            (gt9_rxresetdone_i), // output wire gt9_rxresetdone_i
        //------------------- TX Initialization and Reset Ports --------------------
        .gt9_gttxreset_in               (gt9_gttxreset_i), // input wire gt9_gttxreset_i
        .gt9_txuserrdy_in               (gt9_txuserrdy_i), // input wire gt9_txuserrdy_i
        //-------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        .gt9_txchardispmode_in          (gt9_txchardispmode_in), // input wire [3:0] gt9_txchardispmode_in
        .gt9_txchardispval_in           (gt9_txchardispval_in), // input wire [3:0] gt9_txchardispval_in
        //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
        .gt9_txusrclk_in                (gt9_txusrclk_in), // input wire gt9_txusrclk_in
        .gt9_txusrclk2_in               (gt9_txusrclk2_in), // input wire gt9_txusrclk2_in
        //---------------- Transmit Ports - Pattern Generator Ports ----------------
        .gt9_txprbsforceerr_in          (gt9_txprbsforceerr_in), // input wire gt9_txprbsforceerr_in
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .gt9_txdata_in                  (gt9_txdata_in), // input wire [31:0] gt9_txdata_in
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .gt9_gthtxn_out                 (gt9_gthtxn_out), // output wire gt9_gthtxn_out
        .gt9_gthtxp_out                 (gt9_gthtxp_out), // output wire gt9_gthtxp_out
        //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        .gt9_txoutclk_out               (gt9_txoutclk_i), // output wire gt9_txoutclk_i
        .gt9_txoutclkfabric_out         (gt9_txoutclkfabric_out), // output wire gt9_txoutclkfabric_out
        .gt9_txoutclkpcs_out            (gt9_txoutclkpcs_out), // output wire gt9_txoutclkpcs_out
        //----------- Transmit Ports - TX Initialization and Reset Ports -----------
        .gt9_txresetdone_out            (gt9_txresetdone_i), // output wire gt9_txresetdone_i
        //---------------- Transmit Ports - pattern Generator Ports ----------------
        .gt9_txprbssel_in               (gt9_txprbssel_in), // input wire [2:0] gt9_txprbssel_in
        //--------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        .gt9_txcharisk_in               (gt9_txcharisk_in), // input wire [3:0] gt9_txcharisk_in




    //____________________________COMMON PORTS________________________________
        .gt0_qplloutclk_in              (gt0_qplloutclk_in),
        .gt0_qplloutrefclk_in           (gt0_qplloutrefclk_in),


    //____________________________COMMON PORTS________________________________
        .gt1_qplloutclk_in              (gt1_qplloutclk_in),
        .gt1_qplloutrefclk_in           (gt1_qplloutrefclk_in),


    //____________________________COMMON PORTS________________________________
        .gt2_qplloutclk_in              (gt2_qplloutclk_in),
        .gt2_qplloutrefclk_in           (gt2_qplloutrefclk_in)

    );




assign  gt0_txresetdone_out                  =  gt0_txresetdone_i;
assign  gt0_rxresetdone_out                  =  gt0_rxresetdone_i;
assign  gt0_txoutclk_out                     =  gt0_txoutclk_i;
assign  gt1_txresetdone_out                  =  gt1_txresetdone_i;
assign  gt1_rxresetdone_out                  =  gt1_rxresetdone_i;
assign  gt1_txoutclk_out                     =  gt1_txoutclk_i;
assign  gt3_txresetdone_out                  =  gt3_txresetdone_i;
assign  gt3_rxresetdone_out                  =  gt3_rxresetdone_i;
assign  gt3_txoutclk_out                     =  gt3_txoutclk_i;
assign  gt4_txresetdone_out                  =  gt4_txresetdone_i;
assign  gt4_rxresetdone_out                  =  gt4_rxresetdone_i;
assign  gt4_txoutclk_out                     =  gt4_txoutclk_i;
assign  gt5_txresetdone_out                  =  gt5_txresetdone_i;
assign  gt5_rxresetdone_out                  =  gt5_rxresetdone_i;
assign  gt5_txoutclk_out                     =  gt5_txoutclk_i;
assign  gt7_txresetdone_out                  =  gt7_txresetdone_i;
assign  gt7_rxresetdone_out                  =  gt7_rxresetdone_i;
assign  gt7_txoutclk_out                     =  gt7_txoutclk_i;
assign  gt8_txresetdone_out                  =  gt8_txresetdone_i;
assign  gt8_rxresetdone_out                  =  gt8_rxresetdone_i;
assign  gt8_txoutclk_out                     =  gt8_txoutclk_i;
assign  gt9_txresetdone_out                  =  gt9_txresetdone_i;
assign  gt9_rxresetdone_out                  =  gt9_rxresetdone_i;
assign  gt9_txoutclk_out                     =  gt9_txoutclk_i;
assign  gt0_qpllreset_out                    =  gt0_qpllreset_t;
assign  gt1_qpllreset_out                    =  gt1_qpllreset_t;
assign  gt2_qpllreset_out                    =  gt2_qpllreset_t;

//Assign the outputs from unused (absent) channels to some active signals in case they are ORed together at a higher level
assign  gt2_txresetdone_out                  =  gt0_txresetdone_i;
assign  gt2_rxresetdone_out                  =  gt0_rxresetdone_i;
assign  gt2_txoutclk_out                     =  gt0_txoutclk_i;
assign  gt6_txresetdone_out                  =  gt0_txresetdone_i;
assign  gt6_rxresetdone_out                  =  gt0_rxresetdone_i;
assign  gt6_txoutclk_out                     =  gt0_txoutclk_i;

generate
if (EXAMPLE_USE_CHIPSCOPE == 1) 
begin : chipscope
assign  gt0_gttxreset_i                      =  gt0_gttxreset_in || gt0_gttxreset_t;
assign  gt0_gtrxreset_i                      =  gt0_gtrxreset_in || gt0_gtrxreset_t;
assign  gt0_txuserrdy_i                      =  gt0_txuserrdy_in || gt0_txuserrdy_t;
assign  gt0_rxuserrdy_i                      =  gt0_rxuserrdy_in || gt0_rxuserrdy_t;
assign  gt1_gttxreset_i                      =  gt1_gttxreset_in || gt1_gttxreset_t;
assign  gt1_gtrxreset_i                      =  gt1_gtrxreset_in || gt1_gtrxreset_t;
assign  gt1_txuserrdy_i                      =  gt1_txuserrdy_in || gt1_txuserrdy_t;
assign  gt1_rxuserrdy_i                      =  gt1_rxuserrdy_in || gt1_rxuserrdy_t;
assign  gt2_gttxreset_i                      =  gt2_gttxreset_in || gt2_gttxreset_t;
assign  gt2_gtrxreset_i                      =  gt2_gtrxreset_in || gt2_gtrxreset_t;
assign  gt2_txuserrdy_i                      =  gt2_txuserrdy_in || gt2_txuserrdy_t;
assign  gt2_rxuserrdy_i                      =  gt2_rxuserrdy_in || gt2_rxuserrdy_t;
assign  gt3_gttxreset_i                      =  gt3_gttxreset_in || gt3_gttxreset_t;
assign  gt3_gtrxreset_i                      =  gt3_gtrxreset_in || gt3_gtrxreset_t;
assign  gt3_txuserrdy_i                      =  gt3_txuserrdy_in || gt3_txuserrdy_t;
assign  gt3_rxuserrdy_i                      =  gt3_rxuserrdy_in || gt3_rxuserrdy_t;
assign  gt4_gttxreset_i                      =  gt4_gttxreset_in || gt4_gttxreset_t;
assign  gt4_gtrxreset_i                      =  gt4_gtrxreset_in || gt4_gtrxreset_t;
assign  gt4_txuserrdy_i                      =  gt4_txuserrdy_in || gt4_txuserrdy_t;
assign  gt4_rxuserrdy_i                      =  gt4_rxuserrdy_in || gt4_rxuserrdy_t;
assign  gt5_gttxreset_i                      =  gt5_gttxreset_in || gt5_gttxreset_t;
assign  gt5_gtrxreset_i                      =  gt5_gtrxreset_in || gt5_gtrxreset_t;
assign  gt5_txuserrdy_i                      =  gt5_txuserrdy_in || gt5_txuserrdy_t;
assign  gt5_rxuserrdy_i                      =  gt5_rxuserrdy_in || gt5_rxuserrdy_t;
assign  gt6_gttxreset_i                      =  gt6_gttxreset_in || gt6_gttxreset_t;
assign  gt6_gtrxreset_i                      =  gt6_gtrxreset_in || gt6_gtrxreset_t;
assign  gt6_txuserrdy_i                      =  gt6_txuserrdy_in || gt6_txuserrdy_t;
assign  gt6_rxuserrdy_i                      =  gt6_rxuserrdy_in || gt6_rxuserrdy_t;
assign  gt7_gttxreset_i                      =  gt7_gttxreset_in || gt7_gttxreset_t;
assign  gt7_gtrxreset_i                      =  gt7_gtrxreset_in || gt7_gtrxreset_t;
assign  gt7_txuserrdy_i                      =  gt7_txuserrdy_in || gt7_txuserrdy_t;
assign  gt7_rxuserrdy_i                      =  gt7_rxuserrdy_in || gt7_rxuserrdy_t;
assign  gt8_gttxreset_i                      =  gt8_gttxreset_in || gt8_gttxreset_t;
assign  gt8_gtrxreset_i                      =  gt8_gtrxreset_in || gt8_gtrxreset_t;
assign  gt8_txuserrdy_i                      =  gt8_txuserrdy_in || gt8_txuserrdy_t;
assign  gt8_rxuserrdy_i                      =  gt8_rxuserrdy_in || gt8_rxuserrdy_t;
assign  gt9_gttxreset_i                      =  gt9_gttxreset_in || gt9_gttxreset_t;
assign  gt9_gtrxreset_i                      =  gt9_gtrxreset_in || gt9_gtrxreset_t;
assign  gt9_txuserrdy_i                      =  gt9_txuserrdy_in || gt9_txuserrdy_t;
assign  gt9_rxuserrdy_i                      =  gt9_rxuserrdy_in || gt9_rxuserrdy_t;
end
endgenerate 

generate
if (EXAMPLE_USE_CHIPSCOPE == 0) 
begin : no_chipscope
assign  gt0_gttxreset_i                      =  gt0_gttxreset_t;
assign  gt0_gtrxreset_i                      =  gt0_gtrxreset_t;
assign  gt0_txuserrdy_i                      =  gt0_txuserrdy_t;
assign  gt0_rxuserrdy_i                      =  gt0_rxuserrdy_t;
assign  gt1_gttxreset_i                      =  gt1_gttxreset_t;
assign  gt1_gtrxreset_i                      =  gt1_gtrxreset_t;
assign  gt1_txuserrdy_i                      =  gt1_txuserrdy_t;
assign  gt1_rxuserrdy_i                      =  gt1_rxuserrdy_t;
assign  gt2_gttxreset_i                      =  gt2_gttxreset_t;
assign  gt2_gtrxreset_i                      =  gt2_gtrxreset_t;
assign  gt2_txuserrdy_i                      =  gt2_txuserrdy_t;
assign  gt2_rxuserrdy_i                      =  gt2_rxuserrdy_t;
assign  gt3_gttxreset_i                      =  gt3_gttxreset_t;
assign  gt3_gtrxreset_i                      =  gt3_gtrxreset_t;
assign  gt3_txuserrdy_i                      =  gt3_txuserrdy_t;
assign  gt3_rxuserrdy_i                      =  gt3_rxuserrdy_t;
assign  gt4_gttxreset_i                      =  gt4_gttxreset_t;
assign  gt4_gtrxreset_i                      =  gt4_gtrxreset_t;
assign  gt4_txuserrdy_i                      =  gt4_txuserrdy_t;
assign  gt4_rxuserrdy_i                      =  gt4_rxuserrdy_t;
assign  gt5_gttxreset_i                      =  gt5_gttxreset_t;
assign  gt5_gtrxreset_i                      =  gt5_gtrxreset_t;
assign  gt5_txuserrdy_i                      =  gt5_txuserrdy_t;
assign  gt5_rxuserrdy_i                      =  gt5_rxuserrdy_t;
assign  gt6_gttxreset_i                      =  gt6_gttxreset_t;
assign  gt6_gtrxreset_i                      =  gt6_gtrxreset_t;
assign  gt6_txuserrdy_i                      =  gt6_txuserrdy_t;
assign  gt6_rxuserrdy_i                      =  gt6_rxuserrdy_t;
assign  gt7_gttxreset_i                      =  gt7_gttxreset_t;
assign  gt7_gtrxreset_i                      =  gt7_gtrxreset_t;
assign  gt7_txuserrdy_i                      =  gt7_txuserrdy_t;
assign  gt7_rxuserrdy_i                      =  gt7_rxuserrdy_t;
assign  gt8_gttxreset_i                      =  gt8_gttxreset_t;
assign  gt8_gtrxreset_i                      =  gt8_gtrxreset_t;
assign  gt8_txuserrdy_i                      =  gt8_txuserrdy_t;
assign  gt8_rxuserrdy_i                      =  gt8_rxuserrdy_t;
assign  gt9_gttxreset_i                      =  gt9_gttxreset_t;
assign  gt9_gtrxreset_i                      =  gt9_gtrxreset_t;
assign  gt9_txuserrdy_i                      =  gt9_txuserrdy_t;
assign  gt9_rxuserrdy_i                      =  gt9_rxuserrdy_t;
end
endgenerate 


gtwizard_0_TX_STARTUP_FSM #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),           // Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("TRUE"),                        // the TX and RX Reset FSMs must 
           .RX_QPLL_USED             ("TRUE"),                        // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")               // Decision if a manual phase-alignment is necessary or the automatic 
                                                                     // is enough. For single-lane applications the automatic alignment is 
                                                                     // sufficient              
             ) 
gt0_txresetfsm_i      
            ( 
        .STABLE_CLOCK                   (sysclk_in),
        .TXUSERCLK                      (gt0_txusrclk_in),
        .SOFT_RESET                     (soft_reset_in),
        .QPLLREFCLKLOST                 (gt1_qpllrefclklost_in),
        .CPLLREFCLKLOST                 (tied_to_ground_i),
        .QPLLLOCK                       (gt1_qplllock_in),
        .CPLLLOCK                       (tied_to_vcc_i),
        .TXRESETDONE                    (gt0_txresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .GTTXRESET                      (gt0_gttxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (gt0_qpllreset_t),
        .CPLL_RESET                     (),
        .TX_FSM_RESET_DONE              (gt0_tx_fsm_reset_done_out),
        .TXUSERRDY                      (gt0_txuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RETRY_COUNTER                  ()
           );


gtwizard_0_TX_STARTUP_FSM #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),           // Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("TRUE"),                        // the TX and RX Reset FSMs must 
           .RX_QPLL_USED             ("TRUE"),                        // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")               // Decision if a manual phase-alignment is necessary or the automatic 
                                                                     // is enough. For single-lane applications the automatic alignment is 
                                                                     // sufficient              
             ) 
gt1_txresetfsm_i      
            ( 
        .STABLE_CLOCK                   (sysclk_in),
        .TXUSERCLK                      (gt1_txusrclk_in),
        .SOFT_RESET                     (soft_reset_in),
        .QPLLREFCLKLOST                 (gt2_qpllrefclklost_in),
        .CPLLREFCLKLOST                 (tied_to_ground_i),
        .QPLLLOCK                       (gt2_qplllock_in),
        .CPLLLOCK                       (tied_to_vcc_i),
        .TXRESETDONE                    (gt1_txresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .GTTXRESET                      (gt1_gttxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .TX_FSM_RESET_DONE              (gt1_tx_fsm_reset_done_out),
        .TXUSERRDY                      (gt1_txuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RETRY_COUNTER                  ()
           );

/*
gtwizard_0_TX_STARTUP_FSM #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),           // Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("TRUE"),                        // the TX and RX Reset FSMs must 
           .RX_QPLL_USED             ("TRUE"),                        // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")               // Decision if a manual phase-alignment is necessary or the automatic 
                                                                     // is enough. For single-lane applications the automatic alignment is 
                                                                     // sufficient              
             ) 
gt2_txresetfsm_i      
            ( 
        .STABLE_CLOCK                   (sysclk_in),
        .TXUSERCLK                      (gt2_txusrclk_in),
        .SOFT_RESET                     (soft_reset_in),
        .QPLLREFCLKLOST                 (gt1_qpllrefclklost_in),
        .CPLLREFCLKLOST                 (tied_to_ground_i),
        .QPLLLOCK                       (gt1_qplllock_in),
        .CPLLLOCK                       (tied_to_vcc_i),
        .TXRESETDONE                    (gt2_txresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .GTTXRESET                      (gt2_gttxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (gt1_qpllreset_t),
        .CPLL_RESET                     (),
        .TX_FSM_RESET_DONE              (gt2_tx_fsm_reset_done_out),
        .TXUSERRDY                      (gt2_txuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RETRY_COUNTER                  ()
           );

*/
assign gt2_gttxreset_t = 1'b0;
assign gt2_txuserrdy_t = 1'b1;
assign gt2_tx_fsm_reset_done_out = 1'b1;

gtwizard_0_TX_STARTUP_FSM #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),           // Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("TRUE"),                        // the TX and RX Reset FSMs must 
           .RX_QPLL_USED             ("TRUE"),                        // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")               // Decision if a manual phase-alignment is necessary or the automatic 
                                                                     // is enough. For single-lane applications the automatic alignment is 
                                                                     // sufficient              
             ) 
gt3_txresetfsm_i      
            ( 
        .STABLE_CLOCK                   (sysclk_in),
        .TXUSERCLK                      (gt3_txusrclk_in),
        .SOFT_RESET                     (soft_reset_in),
        .QPLLREFCLKLOST                 (gt2_qpllrefclklost_in),
        .CPLLREFCLKLOST                 (tied_to_ground_i),
        .QPLLLOCK                       (gt2_qplllock_in),
        .CPLLLOCK                       (tied_to_vcc_i),
        .TXRESETDONE                    (gt3_txresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .GTTXRESET                      (gt3_gttxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .TX_FSM_RESET_DONE              (gt3_tx_fsm_reset_done_out),
        .TXUSERRDY                      (gt3_txuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RETRY_COUNTER                  ()
           );


gtwizard_0_TX_STARTUP_FSM #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),           // Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("TRUE"),                        // the TX and RX Reset FSMs must 
           .RX_QPLL_USED             ("TRUE"),                        // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")               // Decision if a manual phase-alignment is necessary or the automatic 
                                                                     // is enough. For single-lane applications the automatic alignment is 
                                                                     // sufficient              
             ) 
gt4_txresetfsm_i      
            ( 
        .STABLE_CLOCK                   (sysclk_in),
        .TXUSERCLK                      (gt4_txusrclk_in),
        .SOFT_RESET                     (soft_reset_in),
        .QPLLREFCLKLOST                 (gt1_qpllrefclklost_in),
        .CPLLREFCLKLOST                 (tied_to_ground_i),
        .QPLLLOCK                       (gt1_qplllock_in),
        .CPLLLOCK                       (tied_to_vcc_i),
        .TXRESETDONE                    (gt4_txresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .GTTXRESET                      (gt4_gttxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .TX_FSM_RESET_DONE              (gt4_tx_fsm_reset_done_out),
        .TXUSERRDY                      (gt4_txuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RETRY_COUNTER                  ()
           );


gtwizard_0_TX_STARTUP_FSM #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),           // Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("TRUE"),                        // the TX and RX Reset FSMs must 
           .RX_QPLL_USED             ("TRUE"),                        // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")               // Decision if a manual phase-alignment is necessary or the automatic 
                                                                     // is enough. For single-lane applications the automatic alignment is 
                                                                     // sufficient              
             ) 
gt5_txresetfsm_i      
            ( 
        .STABLE_CLOCK                   (sysclk_in),
        .TXUSERCLK                      (gt5_txusrclk_in),
        .SOFT_RESET                     (soft_reset_in),
        .QPLLREFCLKLOST                 (gt2_qpllrefclklost_in),
        .CPLLREFCLKLOST                 (tied_to_ground_i),
        .QPLLLOCK                       (gt2_qplllock_in),
        .CPLLLOCK                       (tied_to_vcc_i),
        .TXRESETDONE                    (gt5_txresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .GTTXRESET                      (gt5_gttxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .TX_FSM_RESET_DONE              (gt5_tx_fsm_reset_done_out),
        .TXUSERRDY                      (gt5_txuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RETRY_COUNTER                  ()
           );

/*
gtwizard_0_TX_STARTUP_FSM #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),           // Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("TRUE"),                        // the TX and RX Reset FSMs must 
           .RX_QPLL_USED             ("TRUE"),                        // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")               // Decision if a manual phase-alignment is necessary or the automatic 
                                                                     // is enough. For single-lane applications the automatic alignment is 
                                                                     // sufficient              
             ) 
gt6_txresetfsm_i      
            ( 
        .STABLE_CLOCK                   (sysclk_in),
        .TXUSERCLK                      (gt6_txusrclk_in),
        .SOFT_RESET                     (soft_reset_in),
        .QPLLREFCLKLOST                 (gt2_qpllrefclklost_in),
        .CPLLREFCLKLOST                 (tied_to_ground_i),
        .QPLLLOCK                       (gt2_qplllock_in),
        .CPLLLOCK                       (tied_to_vcc_i),
        .TXRESETDONE                    (gt6_txresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .GTTXRESET                      (gt6_gttxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (gt2_qpllreset_t),
        .CPLL_RESET                     (),
        .TX_FSM_RESET_DONE              (gt6_tx_fsm_reset_done_out),
        .TXUSERRDY                      (gt6_txuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RETRY_COUNTER                  ()
           );
*/
assign gt6_gttxreset_t = 1'b0;
assign gt6_txuserrdy_t = 1'b1;
assign gt6_tx_fsm_reset_done_out = 1'b1;

gtwizard_0_TX_STARTUP_FSM #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),           // Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("TRUE"),                        // the TX and RX Reset FSMs must 
           .RX_QPLL_USED             ("TRUE"),                        // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")               // Decision if a manual phase-alignment is necessary or the automatic 
                                                                     // is enough. For single-lane applications the automatic alignment is 
                                                                     // sufficient              
             ) 
gt7_txresetfsm_i      
            ( 
        .STABLE_CLOCK                   (sysclk_in),
        .TXUSERCLK                      (gt7_txusrclk_in),
        .SOFT_RESET                     (soft_reset_in),
        .QPLLREFCLKLOST                 (gt2_qpllrefclklost_in),
        .CPLLREFCLKLOST                 (tied_to_ground_i),
        .QPLLLOCK                       (gt2_qplllock_in),
        .CPLLLOCK                       (tied_to_vcc_i),
        .TXRESETDONE                    (gt7_txresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .GTTXRESET                      (gt7_gttxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .TX_FSM_RESET_DONE              (gt7_tx_fsm_reset_done_out),
        .TXUSERRDY                      (gt7_txuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RETRY_COUNTER                  ()
           );


gtwizard_0_TX_STARTUP_FSM #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),           // Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("TRUE"),                        // the TX and RX Reset FSMs must 
           .RX_QPLL_USED             ("TRUE"),                        // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")               // Decision if a manual phase-alignment is necessary or the automatic 
                                                                     // is enough. For single-lane applications the automatic alignment is 
                                                                     // sufficient              
             ) 
gt8_txresetfsm_i      
            ( 
        .STABLE_CLOCK                   (sysclk_in),
        .TXUSERCLK                      (gt8_txusrclk_in),
        .SOFT_RESET                     (soft_reset_in),
        .QPLLREFCLKLOST                 (gt1_qpllrefclklost_in),
        .CPLLREFCLKLOST                 (tied_to_ground_i),
        .QPLLLOCK                       (gt1_qplllock_in),
        .CPLLLOCK                       (tied_to_vcc_i),
        .TXRESETDONE                    (gt8_txresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .GTTXRESET                      (gt8_gttxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .TX_FSM_RESET_DONE              (gt8_tx_fsm_reset_done_out),
        .TXUSERRDY                      (gt8_txuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RETRY_COUNTER                  ()
           );


gtwizard_0_TX_STARTUP_FSM #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),           // Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("TRUE"),                        // the TX and RX Reset FSMs must 
           .RX_QPLL_USED             ("TRUE"),                        // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")               // Decision if a manual phase-alignment is necessary or the automatic 
                                                                     // is enough. For single-lane applications the automatic alignment is 
                                                                     // sufficient              
             ) 
gt9_txresetfsm_i      
            ( 
        .STABLE_CLOCK                   (sysclk_in),
        .TXUSERCLK                      (gt9_txusrclk_in),
        .SOFT_RESET                     (soft_reset_in),
        .QPLLREFCLKLOST                 (gt1_qpllrefclklost_in),
        .CPLLREFCLKLOST                 (tied_to_ground_i),
        .QPLLLOCK                       (gt1_qplllock_in),
        .CPLLLOCK                       (tied_to_vcc_i),
        .TXRESETDONE                    (gt9_txresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .GTTXRESET                      (gt9_gttxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .TX_FSM_RESET_DONE              (gt9_tx_fsm_reset_done_out),
        .TXUSERRDY                      (gt9_txuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RETRY_COUNTER                  ()
           );






gtwizard_0_RX_STARTUP_FSM  #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .EQ_MODE                  ("DFE"),                   //Rx Equalization Mode - Set to DFE or LPM
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),              //Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("TRUE"),                           // the TX and RX Reset FSMs must 
           .RX_QPLL_USED             ("TRUE"),                           // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")                 // Decision if a manual phase-alignment is necessary or the automatic 
                                                                         // is enough. For single-lane applications the automatic alignment is 
                                                                         // sufficient              
             )     
gt0_rxresetfsm_i
             ( 
        .STABLE_CLOCK                   (sysclk_in),
        .RXUSERCLK                      (gt0_rxusrclk_in),
        .SOFT_RESET                     (soft_reset_in),
        .RXPMARESETDONE                 (gt0_rxpmaresetdone_i),
        .RXOUTCLK                       (gt0_rxusrclk_in),
        .TXPMARESETDONE                 (gt0_txpmaresetdone_i),
        .TXOUTCLK                       (gt0_txusrclk_in),
        .DONT_RESET_ON_DATA_ERROR       (dont_reset_on_data_error_in),
        .QPLLREFCLKLOST                 (gt1_qpllrefclklost_in),
        .CPLLREFCLKLOST                 (tied_to_ground_i),
        .QPLLLOCK                       (gt1_qplllock_in),
        .CPLLLOCK                       (tied_to_vcc_i),
        .RXRESETDONE                    (gt0_rxresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .RECCLK_STABLE                  (gt0_recclk_stable_i),
        .RECCLK_MONITOR_RESTART         (tied_to_ground_i),
        .DATA_VALID                     (gt0_data_valid_in),
        .TXUSERRDY                      (gt0_txuserrdy_i),
        .GTRXRESET                      (gt0_gtrxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .RX_FSM_RESET_DONE              (gt0_rx_fsm_reset_done_out),
        .RXUSERRDY                      (gt0_rxuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RXDFEAGCHOLD                   (gt0_rxdfeagchold_i),
        .RXDFELFHOLD                    (gt0_rxdfelfhold_i),
        .RXLPMLFHOLD                    (gt0_rxlpmlfhold_i),
        .RXLPMHFHOLD                    (gt0_rxlpmhfhold_i),
        .RETRY_COUNTER                  ()
           );

gtwizard_0_RX_STARTUP_FSM  #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .EQ_MODE                  ("DFE"),                   //Rx Equalization Mode - Set to DFE or LPM
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),              //Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("TRUE"),                           // the TX and RX Reset FSMs must 
           .RX_QPLL_USED             ("TRUE"),                           // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")                 // Decision if a manual phase-alignment is necessary or the automatic 
                                                                         // is enough. For single-lane applications the automatic alignment is 
                                                                         // sufficient              
             )     
gt1_rxresetfsm_i
             ( 
        .STABLE_CLOCK                   (sysclk_in),
        .RXUSERCLK                      (gt1_rxusrclk_in),
        .SOFT_RESET                     (soft_reset_in),
        .RXPMARESETDONE                 (gt0_rxpmaresetdone_i),
        .RXOUTCLK                       (gt1_rxusrclk_in),
        .TXPMARESETDONE                 (gt1_txpmaresetdone_i),
        .TXOUTCLK                       (gt1_txusrclk_in),
        .DONT_RESET_ON_DATA_ERROR       (dont_reset_on_data_error_in),
        .QPLLREFCLKLOST                 (gt2_qpllrefclklost_in),
        .CPLLREFCLKLOST                 (tied_to_ground_i),
        .QPLLLOCK                       (gt2_qplllock_in),
        .CPLLLOCK                       (tied_to_vcc_i),
        .RXRESETDONE                    (gt1_rxresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .RECCLK_STABLE                  (gt0_recclk_stable_i),
        .RECCLK_MONITOR_RESTART         (tied_to_ground_i),
        .DATA_VALID                     (gt1_data_valid_in),
        .TXUSERRDY                      (gt1_txuserrdy_i),
        .GTRXRESET                      (gt1_gtrxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .RX_FSM_RESET_DONE              (gt1_rx_fsm_reset_done_out),
        .RXUSERRDY                      (gt1_rxuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RXDFEAGCHOLD                   (gt1_rxdfeagchold_i),
        .RXDFELFHOLD                    (gt1_rxdfelfhold_i),
        .RXLPMLFHOLD                    (gt1_rxlpmlfhold_i),
        .RXLPMHFHOLD                    (gt1_rxlpmhfhold_i),
        .RETRY_COUNTER                  ()
           );
/*
gtwizard_0_RX_STARTUP_FSM  #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .EQ_MODE                  ("DFE"),                   //Rx Equalization Mode - Set to DFE or LPM
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),              //Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("TRUE"),                           // the TX and RX Reset FSMs must 
           .RX_QPLL_USED             ("TRUE"),                           // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")                 // Decision if a manual phase-alignment is necessary or the automatic 
                                                                         // is enough. For single-lane applications the automatic alignment is 
                                                                         // sufficient              
             )     
gt2_rxresetfsm_i
             ( 
        .STABLE_CLOCK                   (sysclk_in),
        .RXUSERCLK                      (gt2_rxusrclk_in),
        .SOFT_RESET                     (soft_reset_in),
        .RXPMARESETDONE                 (gt0_rxpmaresetdone_i),
        .RXOUTCLK                       (gt2_rxusrclk_in),
        .TXPMARESETDONE                 (gt2_txpmaresetdone_i),
        .TXOUTCLK                       (gt2_txusrclk_in),
        .DONT_RESET_ON_DATA_ERROR       (dont_reset_on_data_error_in),
        .QPLLREFCLKLOST                 (gt1_qpllrefclklost_in),
        .CPLLREFCLKLOST                 (tied_to_ground_i),
        .QPLLLOCK                       (gt1_qplllock_in),
        .CPLLLOCK                       (tied_to_vcc_i),
        .RXRESETDONE                    (gt2_rxresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .RECCLK_STABLE                  (gt0_recclk_stable_i),
        .RECCLK_MONITOR_RESTART         (tied_to_ground_i),
        .DATA_VALID                     (gt2_data_valid_in),
        .TXUSERRDY                      (gt2_txuserrdy_i),
        .GTRXRESET                      (gt2_gtrxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .RX_FSM_RESET_DONE              (gt2_rx_fsm_reset_done_out),
        .RXUSERRDY                      (gt2_rxuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RXDFEAGCHOLD                   (gt2_rxdfeagchold_i),
        .RXDFELFHOLD                    (gt2_rxdfelfhold_i),
        .RXLPMLFHOLD                    (gt2_rxlpmlfhold_i),
        .RXLPMHFHOLD                    (gt2_rxlpmhfhold_i),
        .RETRY_COUNTER                  ()
           );
*/
assign gt2_gtrxreset_t = 1'b0;
assign gt2_rx_fsm_reset_done_out = 1'b1;
assign gt2_rxuserrdy_t = 1'b1;
assign gt2_rxdfeagchold_i = 1'b0;
assign gt2_rxdfelfhold_i = 1'b0;
assign gt2_rxlpmlfhold_i = 1'b0;
assign gt2_rxlpmhfhold_i = 1'b0;

gtwizard_0_RX_STARTUP_FSM  #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .EQ_MODE                  ("DFE"),                   //Rx Equalization Mode - Set to DFE or LPM
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),              //Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("TRUE"),                           // the TX and RX Reset FSMs must 
           .RX_QPLL_USED             ("TRUE"),                           // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")                 // Decision if a manual phase-alignment is necessary or the automatic 
                                                                         // is enough. For single-lane applications the automatic alignment is 
                                                                         // sufficient              
             )     
gt3_rxresetfsm_i
             ( 
        .STABLE_CLOCK                   (sysclk_in),
        .RXUSERCLK                      (gt3_rxusrclk_in),
        .SOFT_RESET                     (soft_reset_in),
        .RXPMARESETDONE                 (gt0_rxpmaresetdone_i),
        .RXOUTCLK                       (gt3_rxusrclk_in),
        .TXPMARESETDONE                 (gt3_txpmaresetdone_i),
        .TXOUTCLK                       (gt3_txusrclk_in),
        .DONT_RESET_ON_DATA_ERROR       (dont_reset_on_data_error_in),
        .QPLLREFCLKLOST                 (gt2_qpllrefclklost_in),
        .CPLLREFCLKLOST                 (tied_to_ground_i),
        .QPLLLOCK                       (gt2_qplllock_in),
        .CPLLLOCK                       (tied_to_vcc_i),
        .RXRESETDONE                    (gt3_rxresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .RECCLK_STABLE                  (gt0_recclk_stable_i),
        .RECCLK_MONITOR_RESTART         (tied_to_ground_i),
        .DATA_VALID                     (gt3_data_valid_in),
        .TXUSERRDY                      (gt3_txuserrdy_i),
        .GTRXRESET                      (gt3_gtrxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .RX_FSM_RESET_DONE              (gt3_rx_fsm_reset_done_out),
        .RXUSERRDY                      (gt3_rxuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RXDFEAGCHOLD                   (gt3_rxdfeagchold_i),
        .RXDFELFHOLD                    (gt3_rxdfelfhold_i),
        .RXLPMLFHOLD                    (gt3_rxlpmlfhold_i),
        .RXLPMHFHOLD                    (gt3_rxlpmhfhold_i),
        .RETRY_COUNTER                  ()
           );

gtwizard_0_RX_STARTUP_FSM  #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .EQ_MODE                  ("DFE"),                   //Rx Equalization Mode - Set to DFE or LPM
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),              //Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("TRUE"),                           // the TX and RX Reset FSMs must 
           .RX_QPLL_USED             ("TRUE"),                           // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")                 // Decision if a manual phase-alignment is necessary or the automatic 
                                                                         // is enough. For single-lane applications the automatic alignment is 
                                                                         // sufficient              
             )     
gt4_rxresetfsm_i
             ( 
        .STABLE_CLOCK                   (sysclk_in),
        .RXUSERCLK                      (gt4_rxusrclk_in),
        .SOFT_RESET                     (soft_reset_in),
        .RXPMARESETDONE                 (gt0_rxpmaresetdone_i),
        .RXOUTCLK                       (gt4_rxusrclk_in),
        .TXPMARESETDONE                 (gt4_txpmaresetdone_i),
        .TXOUTCLK                       (gt4_txusrclk_in),
        .DONT_RESET_ON_DATA_ERROR       (dont_reset_on_data_error_in),
        .QPLLREFCLKLOST                 (gt1_qpllrefclklost_in),
        .CPLLREFCLKLOST                 (tied_to_ground_i),
        .QPLLLOCK                       (gt1_qplllock_in),
        .CPLLLOCK                       (tied_to_vcc_i),
        .RXRESETDONE                    (gt4_rxresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .RECCLK_STABLE                  (gt0_recclk_stable_i),
        .RECCLK_MONITOR_RESTART         (tied_to_ground_i),
        .DATA_VALID                     (gt4_data_valid_in),
        .TXUSERRDY                      (gt4_txuserrdy_i),
        .GTRXRESET                      (gt4_gtrxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .RX_FSM_RESET_DONE              (gt4_rx_fsm_reset_done_out),
        .RXUSERRDY                      (gt4_rxuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RXDFEAGCHOLD                   (gt4_rxdfeagchold_i),
        .RXDFELFHOLD                    (gt4_rxdfelfhold_i),
        .RXLPMLFHOLD                    (gt4_rxlpmlfhold_i),
        .RXLPMHFHOLD                    (gt4_rxlpmhfhold_i),
        .RETRY_COUNTER                  ()
           );

gtwizard_0_RX_STARTUP_FSM  #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .EQ_MODE                  ("DFE"),                   //Rx Equalization Mode - Set to DFE or LPM
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),              //Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("TRUE"),                           // the TX and RX Reset FSMs must 
           .RX_QPLL_USED             ("TRUE"),                           // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")                 // Decision if a manual phase-alignment is necessary or the automatic 
                                                                         // is enough. For single-lane applications the automatic alignment is 
                                                                         // sufficient              
             )     
gt5_rxresetfsm_i
             ( 
        .STABLE_CLOCK                   (sysclk_in),
        .RXUSERCLK                      (gt5_rxusrclk_in),
        .SOFT_RESET                     (soft_reset_in),
        .RXPMARESETDONE                 (gt0_rxpmaresetdone_i),
        .RXOUTCLK                       (gt5_rxusrclk_in),
        .TXPMARESETDONE                 (gt5_txpmaresetdone_i),
        .TXOUTCLK                       (gt5_txusrclk_in),
        .DONT_RESET_ON_DATA_ERROR       (dont_reset_on_data_error_in),
        .QPLLREFCLKLOST                 (gt2_qpllrefclklost_in),
        .CPLLREFCLKLOST                 (tied_to_ground_i),
        .QPLLLOCK                       (gt2_qplllock_in),
        .CPLLLOCK                       (tied_to_vcc_i),
        .RXRESETDONE                    (gt5_rxresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .RECCLK_STABLE                  (gt0_recclk_stable_i),
        .RECCLK_MONITOR_RESTART         (tied_to_ground_i),
        .DATA_VALID                     (gt5_data_valid_in),
        .TXUSERRDY                      (gt5_txuserrdy_i),
        .GTRXRESET                      (gt5_gtrxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .RX_FSM_RESET_DONE              (gt5_rx_fsm_reset_done_out),
        .RXUSERRDY                      (gt5_rxuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RXDFEAGCHOLD                   (gt5_rxdfeagchold_i),
        .RXDFELFHOLD                    (gt5_rxdfelfhold_i),
        .RXLPMLFHOLD                    (gt5_rxlpmlfhold_i),
        .RXLPMHFHOLD                    (gt5_rxlpmhfhold_i),
        .RETRY_COUNTER                  ()
           );
/*
gtwizard_0_RX_STARTUP_FSM  #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .EQ_MODE                  ("DFE"),                   //Rx Equalization Mode - Set to DFE or LPM
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),              //Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("TRUE"),                           // the TX and RX Reset FSMs must 
           .RX_QPLL_USED             ("TRUE"),                           // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")                 // Decision if a manual phase-alignment is necessary or the automatic 
                                                                         // is enough. For single-lane applications the automatic alignment is 
                                                                         // sufficient              
             )     
gt6_rxresetfsm_i
             ( 
        .STABLE_CLOCK                   (sysclk_in),
        .RXUSERCLK                      (gt6_rxusrclk_in),
        .SOFT_RESET                     (soft_reset_in),
        .RXPMARESETDONE                 (gt0_rxpmaresetdone_i),
        .RXOUTCLK                       (gt6_rxusrclk_in),
        .TXPMARESETDONE                 (gt6_txpmaresetdone_i),
        .TXOUTCLK                       (gt6_txusrclk_in),
        .DONT_RESET_ON_DATA_ERROR       (dont_reset_on_data_error_in),
        .QPLLREFCLKLOST                 (gt2_qpllrefclklost_in),
        .CPLLREFCLKLOST                 (tied_to_ground_i),
        .QPLLLOCK                       (gt2_qplllock_in),
        .CPLLLOCK                       (tied_to_vcc_i),
        .RXRESETDONE                    (gt6_rxresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .RECCLK_STABLE                  (gt0_recclk_stable_i),
        .RECCLK_MONITOR_RESTART         (tied_to_ground_i),
        .DATA_VALID                     (gt6_data_valid_in),
        .TXUSERRDY                      (gt6_txuserrdy_i),
        .GTRXRESET                      (gt6_gtrxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .RX_FSM_RESET_DONE              (gt6_rx_fsm_reset_done_out),
        .RXUSERRDY                      (gt6_rxuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RXDFEAGCHOLD                   (gt6_rxdfeagchold_i),
        .RXDFELFHOLD                    (gt6_rxdfelfhold_i),
        .RXLPMLFHOLD                    (gt6_rxlpmlfhold_i),
        .RXLPMHFHOLD                    (gt6_rxlpmhfhold_i),
        .RETRY_COUNTER                  ()
           );
*/

assign gt6_gtrxreset_t = 1'b0;
assign gt6_rx_fsm_reset_done_out = 1'b1;
assign gt6_rxuserrdy_t = 1'b1;
assign gt6_rxdfeagchold_i = 1'b0;
assign gt6_rxdfelfhold_i = 1'b0;
assign gt6_rxlpmlfhold_i = 1'b0;
assign gt6_rxlpmhfhold_i = 1'b0;

gtwizard_0_RX_STARTUP_FSM  #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .EQ_MODE                  ("DFE"),                   //Rx Equalization Mode - Set to DFE or LPM
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),              //Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("TRUE"),                           // the TX and RX Reset FSMs must 
           .RX_QPLL_USED             ("TRUE"),                           // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")                 // Decision if a manual phase-alignment is necessary or the automatic 
                                                                         // is enough. For single-lane applications the automatic alignment is 
                                                                         // sufficient              
             )     
gt7_rxresetfsm_i
             ( 
        .STABLE_CLOCK                   (sysclk_in),
        .RXUSERCLK                      (gt7_rxusrclk_in),
        .SOFT_RESET                     (soft_reset_in),
        .RXPMARESETDONE                 (gt0_rxpmaresetdone_i),
        .RXOUTCLK                       (gt7_rxusrclk_in),
        .TXPMARESETDONE                 (gt7_txpmaresetdone_i),
        .TXOUTCLK                       (gt7_txusrclk_in),
        .DONT_RESET_ON_DATA_ERROR       (dont_reset_on_data_error_in),
        .QPLLREFCLKLOST                 (gt2_qpllrefclklost_in),
        .CPLLREFCLKLOST                 (tied_to_ground_i),
        .QPLLLOCK                       (gt2_qplllock_in),
        .CPLLLOCK                       (tied_to_vcc_i),
        .RXRESETDONE                    (gt7_rxresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .RECCLK_STABLE                  (gt0_recclk_stable_i),
        .RECCLK_MONITOR_RESTART         (tied_to_ground_i),
        .DATA_VALID                     (gt7_data_valid_in),
        .TXUSERRDY                      (gt7_txuserrdy_i),
        .GTRXRESET                      (gt7_gtrxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .RX_FSM_RESET_DONE              (gt7_rx_fsm_reset_done_out),
        .RXUSERRDY                      (gt7_rxuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RXDFEAGCHOLD                   (gt7_rxdfeagchold_i),
        .RXDFELFHOLD                    (gt7_rxdfelfhold_i),
        .RXLPMLFHOLD                    (gt7_rxlpmlfhold_i),
        .RXLPMHFHOLD                    (gt7_rxlpmhfhold_i),
        .RETRY_COUNTER                  ()
           );

gtwizard_0_RX_STARTUP_FSM  #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .EQ_MODE                  ("DFE"),                   //Rx Equalization Mode - Set to DFE or LPM
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),              //Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("TRUE"),                           // the TX and RX Reset FSMs must 
           .RX_QPLL_USED             ("TRUE"),                           // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")                 // Decision if a manual phase-alignment is necessary or the automatic 
                                                                         // is enough. For single-lane applications the automatic alignment is 
                                                                         // sufficient              
             )     
gt8_rxresetfsm_i
             ( 
        .STABLE_CLOCK                   (sysclk_in),
        .RXUSERCLK                      (gt8_rxusrclk_in),
        .SOFT_RESET                     (soft_reset_in),
        .RXPMARESETDONE                 (gt0_rxpmaresetdone_i),
        .RXOUTCLK                       (gt8_rxusrclk_in),
        .TXPMARESETDONE                 (gt8_txpmaresetdone_i),
        .TXOUTCLK                       (gt8_txusrclk_in),
        .DONT_RESET_ON_DATA_ERROR       (dont_reset_on_data_error_in),
        .QPLLREFCLKLOST                 (gt1_qpllrefclklost_in),
        .CPLLREFCLKLOST                 (tied_to_ground_i),
        .QPLLLOCK                       (gt1_qplllock_in),
        .CPLLLOCK                       (tied_to_vcc_i),
        .RXRESETDONE                    (gt8_rxresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .RECCLK_STABLE                  (gt0_recclk_stable_i),
        .RECCLK_MONITOR_RESTART         (tied_to_ground_i),
        .DATA_VALID                     (gt8_data_valid_in),
        .TXUSERRDY                      (gt8_txuserrdy_i),
        .GTRXRESET                      (gt8_gtrxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .RX_FSM_RESET_DONE              (gt8_rx_fsm_reset_done_out),
        .RXUSERRDY                      (gt8_rxuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RXDFEAGCHOLD                   (gt8_rxdfeagchold_i),
        .RXDFELFHOLD                    (gt8_rxdfelfhold_i),
        .RXLPMLFHOLD                    (gt8_rxlpmlfhold_i),
        .RXLPMHFHOLD                    (gt8_rxlpmhfhold_i),
        .RETRY_COUNTER                  ()
           );

gtwizard_0_RX_STARTUP_FSM  #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .EQ_MODE                  ("DFE"),                   //Rx Equalization Mode - Set to DFE or LPM
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),              //Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("TRUE"),                           // the TX and RX Reset FSMs must 
           .RX_QPLL_USED             ("TRUE"),                           // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")                 // Decision if a manual phase-alignment is necessary or the automatic 
                                                                         // is enough. For single-lane applications the automatic alignment is 
                                                                         // sufficient              
             )     
gt9_rxresetfsm_i
             ( 
        .STABLE_CLOCK                   (sysclk_in),
        .RXUSERCLK                      (gt9_rxusrclk_in),
        .SOFT_RESET                     (soft_reset_in),
        .RXPMARESETDONE                 (gt0_rxpmaresetdone_i),
        .RXOUTCLK                       (gt9_rxusrclk_in),
        .TXPMARESETDONE                 (gt9_txpmaresetdone_i),
        .TXOUTCLK                       (gt9_txusrclk_in),
        .DONT_RESET_ON_DATA_ERROR       (dont_reset_on_data_error_in),
        .QPLLREFCLKLOST                 (gt1_qpllrefclklost_in),
        .CPLLREFCLKLOST                 (tied_to_ground_i),
        .QPLLLOCK                       (gt1_qplllock_in),
        .CPLLLOCK                       (tied_to_vcc_i),
        .RXRESETDONE                    (gt9_rxresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .RECCLK_STABLE                  (gt0_recclk_stable_i),
        .RECCLK_MONITOR_RESTART         (tied_to_ground_i),
        .DATA_VALID                     (gt9_data_valid_in),
        .TXUSERRDY                      (gt9_txuserrdy_i),
        .GTRXRESET                      (gt9_gtrxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .RX_FSM_RESET_DONE              (gt9_rx_fsm_reset_done_out),
        .RXUSERRDY                      (gt9_rxuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RXDFEAGCHOLD                   (gt9_rxdfeagchold_i),
        .RXDFELFHOLD                    (gt9_rxdfelfhold_i),
        .RXLPMLFHOLD                    (gt9_rxlpmlfhold_i),
        .RXLPMHFHOLD                    (gt9_rxlpmhfhold_i),
        .RETRY_COUNTER                  ()
           );

  always @(posedge sysclk_in)
  begin
        if(gt0_gtrxreset_i)
        begin
          gt0_rx_cdrlocked       <= `DLY    1'b0;
          gt0_rx_cdrlock_counter <= `DLY    0;      
        end                
        else if (gt0_rx_cdrlock_counter == WAIT_TIME_CDRLOCK) 
        begin
          gt0_rx_cdrlocked       <= `DLY    1'b1;
          gt0_rx_cdrlock_counter <= `DLY    gt0_rx_cdrlock_counter;
        end
        else
          gt0_rx_cdrlock_counter <= `DLY    gt0_rx_cdrlock_counter + 1;
  end 

  always @(posedge sysclk_in)
  begin
        if(gt1_gtrxreset_i)
        begin
          gt1_rx_cdrlocked       <= `DLY    1'b0;
          gt1_rx_cdrlock_counter <= `DLY    0;      
        end                
        else if (gt1_rx_cdrlock_counter == WAIT_TIME_CDRLOCK) 
        begin
          gt1_rx_cdrlocked       <= `DLY    1'b1;
          gt1_rx_cdrlock_counter <= `DLY    gt1_rx_cdrlock_counter;
        end
        else
          gt1_rx_cdrlock_counter <= `DLY    gt1_rx_cdrlock_counter + 1;
  end 

  always @(posedge sysclk_in)
  begin
        if(gt2_gtrxreset_i)
        begin
          gt2_rx_cdrlocked       <= `DLY    1'b0;
          gt2_rx_cdrlock_counter <= `DLY    0;      
        end                
        else if (gt2_rx_cdrlock_counter == WAIT_TIME_CDRLOCK) 
        begin
          gt2_rx_cdrlocked       <= `DLY    1'b1;
          gt2_rx_cdrlock_counter <= `DLY    gt2_rx_cdrlock_counter;
        end
        else
          gt2_rx_cdrlock_counter <= `DLY    gt2_rx_cdrlock_counter + 1;
  end 

  always @(posedge sysclk_in)
  begin
        if(gt3_gtrxreset_i)
        begin
          gt3_rx_cdrlocked       <= `DLY    1'b0;
          gt3_rx_cdrlock_counter <= `DLY    0;      
        end                
        else if (gt3_rx_cdrlock_counter == WAIT_TIME_CDRLOCK) 
        begin
          gt3_rx_cdrlocked       <= `DLY    1'b1;
          gt3_rx_cdrlock_counter <= `DLY    gt3_rx_cdrlock_counter;
        end
        else
          gt3_rx_cdrlock_counter <= `DLY    gt3_rx_cdrlock_counter + 1;
  end 

  always @(posedge sysclk_in)
  begin
        if(gt4_gtrxreset_i)
        begin
          gt4_rx_cdrlocked       <= `DLY    1'b0;
          gt4_rx_cdrlock_counter <= `DLY    0;      
        end                
        else if (gt4_rx_cdrlock_counter == WAIT_TIME_CDRLOCK) 
        begin
          gt4_rx_cdrlocked       <= `DLY    1'b1;
          gt4_rx_cdrlock_counter <= `DLY    gt4_rx_cdrlock_counter;
        end
        else
          gt4_rx_cdrlock_counter <= `DLY    gt4_rx_cdrlock_counter + 1;
  end 

  always @(posedge sysclk_in)
  begin
        if(gt5_gtrxreset_i)
        begin
          gt5_rx_cdrlocked       <= `DLY    1'b0;
          gt5_rx_cdrlock_counter <= `DLY    0;      
        end                
        else if (gt5_rx_cdrlock_counter == WAIT_TIME_CDRLOCK) 
        begin
          gt5_rx_cdrlocked       <= `DLY    1'b1;
          gt5_rx_cdrlock_counter <= `DLY    gt5_rx_cdrlock_counter;
        end
        else
          gt5_rx_cdrlock_counter <= `DLY    gt5_rx_cdrlock_counter + 1;
  end 

  always @(posedge sysclk_in)
  begin
        if(gt6_gtrxreset_i)
        begin
          gt6_rx_cdrlocked       <= `DLY    1'b0;
          gt6_rx_cdrlock_counter <= `DLY    0;      
        end                
        else if (gt6_rx_cdrlock_counter == WAIT_TIME_CDRLOCK) 
        begin
          gt6_rx_cdrlocked       <= `DLY    1'b1;
          gt6_rx_cdrlock_counter <= `DLY    gt6_rx_cdrlock_counter;
        end
        else
          gt6_rx_cdrlock_counter <= `DLY    gt6_rx_cdrlock_counter + 1;
  end 

  always @(posedge sysclk_in)
  begin
        if(gt7_gtrxreset_i)
        begin
          gt7_rx_cdrlocked       <= `DLY    1'b0;
          gt7_rx_cdrlock_counter <= `DLY    0;      
        end                
        else if (gt7_rx_cdrlock_counter == WAIT_TIME_CDRLOCK) 
        begin
          gt7_rx_cdrlocked       <= `DLY    1'b1;
          gt7_rx_cdrlock_counter <= `DLY    gt7_rx_cdrlock_counter;
        end
        else
          gt7_rx_cdrlock_counter <= `DLY    gt7_rx_cdrlock_counter + 1;
  end 

  always @(posedge sysclk_in)
  begin
        if(gt8_gtrxreset_i)
        begin
          gt8_rx_cdrlocked       <= `DLY    1'b0;
          gt8_rx_cdrlock_counter <= `DLY    0;      
        end                
        else if (gt8_rx_cdrlock_counter == WAIT_TIME_CDRLOCK) 
        begin
          gt8_rx_cdrlocked       <= `DLY    1'b1;
          gt8_rx_cdrlock_counter <= `DLY    gt8_rx_cdrlock_counter;
        end
        else
          gt8_rx_cdrlock_counter <= `DLY    gt8_rx_cdrlock_counter + 1;
  end 

  always @(posedge sysclk_in)
  begin
        if(gt9_gtrxreset_i)
        begin
          gt9_rx_cdrlocked       <= `DLY    1'b0;
          gt9_rx_cdrlock_counter <= `DLY    0;      
        end                
        else if (gt9_rx_cdrlock_counter == WAIT_TIME_CDRLOCK) 
        begin
          gt9_rx_cdrlocked       <= `DLY    1'b1;
          gt9_rx_cdrlock_counter <= `DLY    gt9_rx_cdrlock_counter;
        end
        else
          gt9_rx_cdrlock_counter <= `DLY    gt9_rx_cdrlock_counter + 1;
  end 

assign  gt0_recclk_stable_i                  =  gt0_rx_cdrlocked;
assign  gt1_recclk_stable_i                  =  gt1_rx_cdrlocked;
assign  gt2_recclk_stable_i                  =  gt2_rx_cdrlocked;
assign  gt3_recclk_stable_i                  =  gt3_rx_cdrlocked;
assign  gt4_recclk_stable_i                  =  gt4_rx_cdrlocked;
assign  gt5_recclk_stable_i                  =  gt5_rx_cdrlocked;
assign  gt6_recclk_stable_i                  =  gt6_rx_cdrlocked;
assign  gt7_recclk_stable_i                  =  gt7_rx_cdrlocked;
assign  gt8_recclk_stable_i                  =  gt8_rx_cdrlocked;
assign  gt9_recclk_stable_i                  =  gt9_rx_cdrlocked;







endmodule


